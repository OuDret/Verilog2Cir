.SUBCKT Gaussian VSS VDD clk reset sensor1 sensor2 sensor3 sensor4 sensor5 sensor6 central_value finestra_gaussiana1 finestra_gaussiana2 finestra_gaussiana3 finestra_gaussiana4 finestra_gaussiana5 finestra_gaussiana6
X2560 VSS VDD reset _0016_ INVERTER
X2561 VSS VDD clk _0015_ INVERTER
X2562 VSS VDD sensor4_7_ finestra_gaussiana4_3_ _0287_ NAND2
X2563 VSS VDD _0287_ _0298_ INVERTER
X2564 VSS VDD sensor4_6_ finestra_gaussiana4_4_ _0309_ NAND2
X2565 VSS VDD finestra_gaussiana4_5_ sensor4_5_ _0320_ NAND2
X2566 VSS VDD sensor4_6_ finestra_gaussiana4_5_ _0331_ NAND2
X2567 VSS VDD finestra_gaussiana4_4_ sensor4_5_ _0342_ NAND2
X2568 VSS VDD _0331_ _0342_ _0353_ NOR2
X2569 VSS VDD _0309_ _0320_ _0364_ XOR
X2570 VSS VDD _0298_ _0364_ _0375_ NAND2
X2571 VSS VDD sensor4_7_ finestra_gaussiana4_4_ _0386_ NAND2
X2572 VSS VDD sensor4_7_ finestra_gaussiana4_5_ _0397_ NAND2
X2573 VSS VDD _0309_ _0397_ _0408_ NOR2
X2574 VSS VDD _0331_ _0386_ _0419_ XOR
X2575 VSS VDD _0375_ _0419_ _0430_ XOR
X2576 VSS VDD finestra_gaussiana4_7_ sensor4_4_ _0441_ NAND2
X2577 VSS VDD finestra_gaussiana4_6_ _0353_ _0452_ NAND2
X2578 VSS VDD finestra_gaussiana4_6_ sensor4_5_ _0353_ _0463_ AOI21
X2579 VSS VDD finestra_gaussiana4_6_ _0353_ _0463_ _0474_ AOI21
X2580 VSS VDD finestra_gaussiana4_7_ sensor4_4_ _0474_ _0485_ AOI21
X2581 VSS VDD finestra_gaussiana4_6_ _0353_ _0441_ _0463_ _0496_ AOI211
X2582 VSS VDD finestra_gaussiana4_7_ sensor4_4_ _0474_ _0507_ NAND3
X2583 VSS VDD _0485_ _0496_ _0518_ NOR2
X2584 VSS VDD _0441_ _0474_ _0529_ XOR
X2585 VSS VDD _0430_ _0529_ _0540_ NOR2
X2586 VSS VDD _0298_ _0364_ _0419_ _0540_ _0551_ AOI31
X2587 VSS VDD finestra_gaussiana4_7_ sensor4_5_ _0562_ NAND2
X2588 VSS VDD finestra_gaussiana4_6_ _0408_ _0573_ NAND2
X2589 VSS VDD sensor4_6_ finestra_gaussiana4_6_ _0408_ _0584_ AOI21
X2590 VSS VDD finestra_gaussiana4_6_ _0408_ _0584_ _0595_ AOI21
X2591 VSS VDD _0562_ _0595_ _0606_ XOR
X2592 VSS VDD _0606_ _0617_ INVERTER
X2593 VSS VDD _0397_ _0606_ _0628_ NOR2
X2594 VSS VDD _0397_ _0606_ _0639_ XOR
X2595 VSS VDD _0397_ _0617_ _0650_ XOR
X2596 VSS VDD _0551_ _0650_ _0661_ NOR2
X2597 VSS VDD _0551_ _0639_ _0672_ XOR
X2598 VSS VDD _0441_ _0463_ _0452_ _0683_ OAI21
X2599 VSS VDD _0452_ _0507_ _0672_ _0694_ AOI21
X2600 VSS VDD _0661_ _0694_ _0705_ NOR2
X2601 VSS VDD finestra_gaussiana4_6_ sensor4_7_ _0716_ NAND2
X2602 VSS VDD finestra_gaussiana4_7_ sensor4_6_ _0727_ NAND2
X2603 VSS VDD finestra_gaussiana4_7_ sensor4_7_ _0738_ NAND2
X2604 VSS VDD _0716_ _0727_ _0749_ XOR
X2605 VSS VDD _0628_ _0749_ _0760_ NAND2
X2606 VSS VDD _0628_ _0749_ _0771_ XOR
X2607 VSS VDD _0562_ _0584_ _0573_ _0782_ OAI21
X2608 VSS VDD _0771_ _0782_ _0793_ NAND2
X2609 VSS VDD _0771_ _0782_ _0804_ XOR
X2610 VSS VDD _0661_ _0694_ _0804_ _0815_ OAI21
X2611 VSS VDD sensor4_5_ finestra_gaussiana4_3_ _0826_ NAND2
X2612 VSS VDD sensor4_7_ finestra_gaussiana4_1_ _0837_ NAND2
X2613 VSS VDD sensor4_5_ finestra_gaussiana4_1_ _0848_ NAND2
X2614 VSS VDD _0287_ _0848_ _0859_ NOR2
X2615 VSS VDD sensor4_6_ _0859_ _0870_ NAND2
X2616 VSS VDD sensor4_6_ finestra_gaussiana4_3_ _0881_ NAND2
X2617 VSS VDD sensor4_6_ finestra_gaussiana4_3_ _0859_ _0892_ AOI21
X2618 VSS VDD _0287_ _0848_ _0881_ _0903_ OAI21
X2619 VSS VDD sensor4_6_ _0859_ _0892_ _0914_ AOI21
X2620 VSS VDD _0870_ _0903_ _0925_ NAND2
X2621 VSS VDD finestra_gaussiana4_5_ sensor4_4_ _0936_ NAND2
X2622 VSS VDD sensor4_7_ finestra_gaussiana4_2_ _0947_ NAND2
X2623 VSS VDD sensor4_5_ finestra_gaussiana4_2_ _0958_ NAND2
X2624 VSS VDD _0386_ _0958_ _0969_ NOR2
X2625 VSS VDD _0342_ _0947_ _0980_ XOR
X2626 VSS VDD _0936_ _0980_ _0991_ XOR
X2627 VSS VDD _0892_ _0991_ _0870_ _1002_ OAI21
X2628 VSS VDD _0298_ _0364_ _1013_ XOR
X2629 VSS VDD _0287_ _0364_ _1024_ XOR
X2630 VSS VDD _1002_ _1024_ _1035_ XOR
X2631 VSS VDD finestra_gaussiana4_7_ sensor4_3_ _1046_ NAND2
X2632 VSS VDD finestra_gaussiana4_6_ sensor4_4_ _1057_ NAND2
X2633 VSS VDD finestra_gaussiana4_5_ sensor4_4_ _0980_ _0969_ _1068_ AOI31
X2634 VSS VDD _1057_ _1068_ _1079_ XOR
X2635 VSS VDD finestra_gaussiana4_7_ sensor4_3_ _1079_ _1090_ NAND3
X2636 VSS VDD _1046_ _1079_ _1101_ XOR
X2637 VSS VDD _1035_ _1101_ _1112_ NOR2
X2638 VSS VDD _1002_ _1013_ _1112_ _1123_ AOI21
X2639 VSS VDD _0430_ _0518_ _1134_ XOR
X2640 VSS VDD _1123_ _1134_ _1145_ NOR2
X2641 VSS VDD _1123_ _1134_ _1156_ XOR
X2642 VSS VDD _1057_ _1068_ _1090_ _1167_ OAI21
X2643 VSS VDD _1156_ _1167_ _1145_ _1178_ AOI21
X2644 VSS VDD _0672_ _0683_ _1189_ XOR
X2645 VSS VDD _1189_ _1200_ INVERTER
X2646 VSS VDD _1178_ _1189_ _1211_ NOR2
X2647 VSS VDD sensor4_7_ finestra_gaussiana4_0_ _1222_ NAND2
X2648 VSS VDD finestra_gaussiana4_3_ sensor4_4_ _1233_ NAND2
X2649 VSS VDD sensor4_4_ finestra_gaussiana4_0_ _1244_ NAND2
X2650 VSS VDD _0287_ _1244_ _1255_ NOR2
X2651 VSS VDD _1222_ _1233_ _1266_ XOR
X2652 VSS VDD sensor4_6_ finestra_gaussiana4_1_ _1277_ NAND2
X2653 VSS VDD sensor4_6_ finestra_gaussiana4_1_ _1266_ _1288_ NAND3
X2654 VSS VDD sensor4_6_ finestra_gaussiana4_1_ _1266_ _1255_ _1299_ AOI31
X2655 VSS VDD _0287_ _1244_ _1288_ _1310_ OAI21
X2656 VSS VDD _0826_ _0837_ _1321_ XOR
X2657 VSS VDD _1310_ _1321_ _1332_ NAND2
X2658 VSS VDD _1299_ _1321_ _1343_ XOR
X2659 VSS VDD finestra_gaussiana4_5_ sensor4_3_ _1354_ NAND2
X2660 VSS VDD finestra_gaussiana4_4_ sensor4_4_ _1365_ NAND2
X2661 VSS VDD sensor4_6_ finestra_gaussiana4_2_ _1376_ NAND2
X2662 VSS VDD sensor4_4_ finestra_gaussiana4_2_ _1387_ NAND2
X2663 VSS VDD _0309_ _1387_ _1398_ NOR2
X2664 VSS VDD _1365_ _1376_ _1409_ XOR
X2665 VSS VDD finestra_gaussiana4_5_ sensor4_3_ _1409_ _1420_ NAND3
X2666 VSS VDD _1354_ _1409_ _1431_ XOR
X2667 VSS VDD _1343_ _1431_ _1332_ _1442_ OAI21
X2668 VSS VDD _0925_ _0991_ _1453_ XOR
X2669 VSS VDD _0914_ _0991_ _1464_ XOR
X2670 VSS VDD _1442_ _1453_ _1475_ NAND2
X2671 VSS VDD _1442_ _1464_ _1486_ XOR
X2672 VSS VDD finestra_gaussiana4_7_ sensor4_2_ _1497_ NAND2
X2673 VSS VDD finestra_gaussiana4_6_ sensor4_3_ _1508_ NAND2
X2674 VSS VDD finestra_gaussiana4_5_ sensor4_3_ _1409_ _1398_ _1519_ AOI31
X2675 VSS VDD _0309_ _1387_ _1420_ _1530_ OAI21
X2676 VSS VDD finestra_gaussiana4_6_ sensor4_3_ _1530_ _1541_ NAND3
X2677 VSS VDD _1508_ _1519_ _1552_ XOR
X2678 VSS VDD finestra_gaussiana4_7_ sensor4_2_ _1552_ _1563_ NAND3
X2679 VSS VDD _1497_ _1552_ _1574_ XOR
X2680 VSS VDD _1486_ _1574_ _1475_ _1585_ OAI21
X2681 VSS VDD _1035_ _1101_ _1596_ XOR
X2682 VSS VDD _1585_ _1596_ _1607_ XOR
X2683 VSS VDD _1607_ _1618_ INVERTER
X2684 VSS VDD _1541_ _1563_ _1629_ NAND2
X2685 VSS VDD _1541_ _1563_ _1618_ _1640_ AOI21
X2686 VSS VDD _1585_ _1596_ _1640_ _1651_ AOI21
X2687 VSS VDD _1651_ _1662_ INVERTER
X2688 VSS VDD _1156_ _1167_ _1673_ XOR
X2689 VSS VDD _1662_ _1673_ _1684_ NAND2
X2690 VSS VDD _1651_ _1673_ _1695_ XOR
X2691 VSS VDD sensor4_6_ finestra_gaussiana4_0_ _1706_ NAND2
X2692 VSS VDD finestra_gaussiana4_3_ sensor4_3_ _1717_ NAND2
X2693 VSS VDD sensor4_3_ finestra_gaussiana4_0_ _1728_ NAND2
X2694 VSS VDD _0881_ _1728_ _1739_ NOR2
X2695 VSS VDD _1706_ _1717_ _1750_ XOR
X2696 VSS VDD sensor4_5_ finestra_gaussiana4_1_ _1750_ _1739_ _1761_ AOI31
X2697 VSS VDD _1266_ _1277_ _1772_ XOR
X2698 VSS VDD _1761_ _1772_ _1783_ XOR
X2699 VSS VDD finestra_gaussiana4_5_ sensor4_2_ _1793_ NAND2
X2700 VSS VDD finestra_gaussiana4_4_ sensor4_3_ _1804_ NAND2
X2701 VSS VDD _0958_ _1804_ _1814_ NAND2
X2702 VSS VDD finestra_gaussiana4_2_ sensor4_3_ _1822_ NAND2
X2703 VSS VDD _0342_ _1822_ _1823_ NOR2
X2704 VSS VDD _0342_ _1822_ _1814_ _1824_ OAI21
X2705 VSS VDD _1793_ _1824_ _1825_ XOR
X2706 VSS VDD _1783_ _1825_ _1826_ NAND2
X2707 VSS VDD _1761_ _1772_ _1826_ _1827_ OAI21
X2708 VSS VDD _1343_ _1431_ _1828_ XOR
X2709 VSS VDD _1827_ _1828_ _1829_ NAND2
X2710 VSS VDD _1827_ _1828_ _1830_ NOR2
X2711 VSS VDD _1827_ _1828_ _1831_ XOR
X2712 VSS VDD finestra_gaussiana4_7_ sensor4_1_ _1832_ NAND2
X2713 VSS VDD finestra_gaussiana4_6_ sensor4_2_ _1833_ NAND2
X2714 VSS VDD finestra_gaussiana4_5_ sensor4_2_ _1814_ _1823_ _1834_ AOI31
X2715 VSS VDD _1833_ _1834_ _1835_ XOR
X2716 VSS VDD finestra_gaussiana4_7_ sensor4_1_ _1835_ _1836_ NAND3
X2717 VSS VDD _1832_ _1835_ _1837_ XOR
X2718 VSS VDD _1830_ _1837_ _1829_ _1838_ OAI21
X2719 VSS VDD _1486_ _1574_ _1839_ XOR
X2720 VSS VDD _1838_ _1839_ _1840_ NAND2
X2721 VSS VDD _1838_ _1839_ _1841_ XOR
X2722 VSS VDD _1833_ _1834_ _1836_ _1842_ OAI21
X2723 VSS VDD _1841_ _1842_ _1843_ NAND2
X2724 VSS VDD _1840_ _1843_ _1844_ NAND2
X2725 VSS VDD _1618_ _1629_ _1845_ XOR
X2726 VSS VDD _1840_ _1843_ _1845_ _1846_ AOI21
X2727 VSS VDD _1844_ _1845_ _1847_ XOR
X2728 VSS VDD sensor4_5_ finestra_gaussiana4_0_ _1848_ NAND2
X2729 VSS VDD finestra_gaussiana4_3_ sensor4_2_ _1849_ NAND2
X2730 VSS VDD finestra_gaussiana4_0_ sensor4_2_ _1850_ NAND2
X2731 VSS VDD _0826_ _1850_ _1851_ NOR2
X2732 VSS VDD _1848_ _1849_ _1852_ XOR
X2733 VSS VDD sensor4_4_ finestra_gaussiana4_1_ _1853_ NAND2
X2734 VSS VDD sensor4_4_ finestra_gaussiana4_1_ _1852_ _1851_ _1854_ AOI31
X2735 VSS VDD _0848_ _1750_ _1855_ XOR
X2736 VSS VDD _1854_ _1855_ _1856_ NOR2
X2737 VSS VDD _1854_ _1855_ _1857_ XOR
X2738 VSS VDD finestra_gaussiana4_5_ sensor4_1_ _1858_ NAND2
X2739 VSS VDD finestra_gaussiana4_4_ sensor4_2_ _1859_ NAND2
X2740 VSS VDD finestra_gaussiana4_2_ sensor4_2_ _1860_ NAND2
X2741 VSS VDD _1387_ _1859_ _1861_ NOR2
X2742 VSS VDD _1387_ _1859_ _1862_ NAND2
X2743 VSS VDD _1387_ _1859_ _1863_ XOR
X2744 VSS VDD _1365_ _1860_ _1862_ _1864_ OAI21
X2745 VSS VDD _1858_ _1864_ _1865_ NOR2
X2746 VSS VDD _1858_ _1864_ _1866_ XOR
X2747 VSS VDD _1858_ _1863_ _1867_ XOR
X2748 VSS VDD _1857_ _1866_ _1868_ NAND2
X2749 VSS VDD _1857_ _1866_ _1856_ _1869_ AOI21
X2750 VSS VDD _1854_ _1855_ _1868_ _1870_ OAI21
X2751 VSS VDD _1783_ _1825_ _1871_ XOR
X2752 VSS VDD _1870_ _1871_ _1872_ NAND2
X2753 VSS VDD _1869_ _1871_ _1873_ XOR
X2754 VSS VDD finestra_gaussiana4_7_ sensor4_0_ _1874_ NAND2
X2755 VSS VDD finestra_gaussiana4_6_ sensor4_1_ _1875_ NAND2
X2756 VSS VDD finestra_gaussiana4_5_ sensor4_1_ _1862_ _1861_ _1876_ AOI31
X2757 VSS VDD _1861_ _1865_ finestra_gaussiana4_6_ sensor4_1_ _1877_ OAI211
X2758 VSS VDD _1875_ _1876_ _1878_ XOR
X2759 VSS VDD finestra_gaussiana4_7_ sensor4_0_ _1878_ _1879_ NAND3
X2760 VSS VDD _1874_ _1878_ _1880_ XOR
X2761 VSS VDD _1873_ _1880_ _1872_ _1881_ OAI21
X2762 VSS VDD _1881_ _1882_ INVERTER
X2763 VSS VDD _1831_ _1837_ _1883_ XOR
X2764 VSS VDD _1882_ _1883_ _1884_ NOR2
X2765 VSS VDD _1881_ _1883_ _1885_ XOR
X2766 VSS VDD _1877_ _1879_ _1886_ NAND2
X2767 VSS VDD _1877_ _1879_ _1885_ _1887_ AOI21
X2768 VSS VDD _1884_ _1887_ _1888_ NOR2
X2769 VSS VDD _1888_ _1889_ INVERTER
X2770 VSS VDD _1841_ _1842_ _1890_ XOR
X2771 VSS VDD _1884_ _1887_ _1890_ _1891_ OAI21
X2772 VSS VDD _1889_ _1890_ _1892_ XOR
X2773 VSS VDD _1888_ _1890_ _1893_ XOR
X2774 VSS VDD finestra_gaussiana4_3_ sensor4_1_ _1894_ NAND2
X2775 VSS VDD finestra_gaussiana4_0_ sensor4_1_ _1895_ NAND2
X2776 VSS VDD _1233_ _1895_ _1896_ NOR2
X2777 VSS VDD _1244_ _1894_ _1897_ XOR
X2778 VSS VDD finestra_gaussiana4_1_ sensor4_3_ _1898_ NAND2
X2779 VSS VDD finestra_gaussiana4_1_ sensor4_3_ _1897_ _1896_ _1899_ AOI31
X2780 VSS VDD _1852_ _1853_ _1900_ XOR
X2781 VSS VDD _1899_ _1900_ _1901_ NOR2
X2782 VSS VDD _1899_ _1900_ _1902_ XOR
X2783 VSS VDD finestra_gaussiana4_5_ sensor4_0_ _1903_ NAND2
X2784 VSS VDD finestra_gaussiana4_4_ sensor4_1_ _1904_ NAND2
X2785 VSS VDD finestra_gaussiana4_2_ sensor4_1_ _1905_ NAND2
X2786 VSS VDD _1804_ _1905_ _1906_ NOR2
X2787 VSS VDD _1822_ _1904_ _1907_ NAND2
X2788 VSS VDD _1804_ _1905_ _1907_ _1908_ OAI21
X2789 VSS VDD _1903_ _1908_ _1909_ XOR
X2790 VSS VDD _1902_ _1909_ _1901_ _1910_ AOI21
X2791 VSS VDD _1857_ _1867_ _1911_ XOR
X2792 VSS VDD _1910_ _1911_ _1912_ XOR
X2793 VSS VDD finestra_gaussiana4_6_ sensor4_0_ _1913_ NAND2
X2794 VSS VDD finestra_gaussiana4_5_ sensor4_0_ _1907_ _1906_ _1914_ AOI31
X2795 VSS VDD _1913_ _1914_ _1915_ NOR2
X2796 VSS VDD _1913_ _1914_ _1916_ XOR
X2797 VSS VDD _1912_ _1916_ _1917_ NAND2
X2798 VSS VDD _1910_ _1911_ _1917_ _1918_ OAI21
X2799 VSS VDD _1873_ _1880_ _1919_ XOR
X2800 VSS VDD _1918_ _1919_ _1920_ NAND2
X2801 VSS VDD _1918_ _1919_ _1921_ XOR
X2802 VSS VDD _1915_ _1921_ _1922_ NAND2
X2803 VSS VDD _1920_ _1922_ _1923_ NAND2
X2804 VSS VDD _1885_ _1886_ _1924_ XOR
X2805 VSS VDD _1920_ _1922_ _1924_ _1925_ AOI21
X2806 VSS VDD _1897_ _1898_ _1926_ XOR
X2807 VSS VDD finestra_gaussiana4_3_ sensor4_0_ _1927_ NAND2
X2808 VSS VDD finestra_gaussiana4_0_ sensor4_0_ _1928_ NAND2
X2809 VSS VDD _1717_ _1928_ _1929_ NOR2
X2810 VSS VDD finestra_gaussiana4_1_ sensor4_2_ _1930_ NAND2
X2811 VSS VDD _1728_ _1927_ _1930_ _1931_ AOI21
X2812 VSS VDD _1929_ _1931_ _1932_ NOR2
X2813 VSS VDD _1926_ _1932_ _1933_ NOR2
X2814 VSS VDD finestra_gaussiana4_4_ sensor4_0_ _1934_ NAND2
X2815 VSS VDD finestra_gaussiana4_2_ sensor4_0_ _1935_ NAND2
X2816 VSS VDD _1859_ _1935_ _1936_ NOR2
X2817 VSS VDD _1860_ _1934_ _1937_ XOR
X2818 VSS VDD _1926_ _1932_ _1938_ XOR
X2819 VSS VDD _1937_ _1938_ _1933_ _1939_ AOI21
X2820 VSS VDD _1939_ _1940_ INVERTER
X2821 VSS VDD _1902_ _1909_ _1941_ XOR
X2822 VSS VDD _1940_ _1941_ _1942_ NAND2
X2823 VSS VDD _1940_ _1941_ _1943_ XOR
X2824 VSS VDD _1939_ _1941_ _1944_ XOR
X2825 VSS VDD _1936_ _1943_ _1945_ NAND2
X2826 VSS VDD _1859_ _1935_ _1942_ _1944_ _1946_ OAI31
X2827 VSS VDD _1912_ _1916_ _1947_ XOR
X2828 VSS VDD _1947_ _1948_ INVERTER
X2829 VSS VDD _1942_ _1945_ _1948_ _1949_ AOI21
X2830 VSS VDD _1946_ _1947_ _1950_ NAND2
X2831 VSS VDD _1915_ _1921_ _1951_ XOR
X2832 VSS VDD _1949_ _1951_ _1952_ NAND2
X2833 VSS VDD _1728_ _1927_ _1953_ XOR
X2834 VSS VDD finestra_gaussiana4_1_ sensor4_1_ _1954_ NAND2
X2835 VSS VDD _1895_ _1930_ _1953_ _1955_ NOR3
X2836 VSS VDD finestra_gaussiana4_0_ sensor4_1_ _1930_ _1956_ AOI21
X2837 VSS VDD finestra_gaussiana4_1_ sensor4_2_ _1895_ _1957_ NAND3
X2838 VSS VDD _1953_ _1957_ _1958_ XOR
X2839 VSS VDD _1953_ _1956_ _1959_ XOR
X2840 VSS VDD _1905_ _1958_ _1960_ NOR2
X2841 VSS VDD finestra_gaussiana4_2_ sensor4_1_ _1959_ _1955_ _1961_ AOI31
X2842 VSS VDD _1937_ _1938_ _1962_ XOR
X2843 VSS VDD _1955_ _1960_ _1962_ _1963_ OAI21
X2844 VSS VDD _1936_ _1943_ _1964_ XOR
X2845 VSS VDD _1936_ _1944_ _1965_ XOR
X2846 VSS VDD _1963_ _1965_ _1966_ NOR2
X2847 VSS VDD _1946_ _1947_ _1967_ XOR
X2848 VSS VDD _1946_ _1948_ _1968_ XOR
X2849 VSS VDD _1966_ _1967_ _1969_ NAND2
X2850 VSS VDD finestra_gaussiana4_1_ sensor4_0_ _1970_ NAND2
X2851 VSS VDD _1928_ _1954_ _1971_ NOR2
X2852 VSS VDD _1850_ _1954_ _1972_ XOR
X2853 VSS VDD _1971_ _1972_ _1973_ NAND2
X2854 VSS VDD _1971_ _1972_ _1974_ NOR2
X2855 VSS VDD _1971_ _1972_ _1975_ XOR
X2856 VSS VDD _1935_ _1974_ _1973_ _1976_ OAI21
X2857 VSS VDD _1905_ _1958_ _1977_ XOR
X2858 VSS VDD _1905_ _1959_ _1978_ XOR
X2859 VSS VDD _1976_ _1977_ _1979_ NAND2
X2860 VSS VDD _1961_ _1962_ _1980_ XOR
X2861 VSS VDD _1979_ _1980_ _1981_ NOR2
X2862 VSS VDD _1964_ _1981_ _1982_ NAND2
X2863 VSS VDD _1966_ _1968_ _1983_ XOR
X2864 VSS VDD _1982_ _1983_ _1969_ _1984_ OAI21
X2865 VSS VDD _1949_ _1951_ _1985_ XOR
X2866 VSS VDD _1950_ _1951_ _1986_ XOR
X2867 VSS VDD _1984_ _1985_ _1987_ NAND2
X2868 VSS VDD _1952_ _1987_ _1988_ NAND2
X2869 VSS VDD _1923_ _1924_ _1989_ XOR
X2870 VSS VDD _1989_ _1990_ INVERTER
X2871 VSS VDD _1952_ _1987_ _1989_ _1991_ AOI21
X2872 VSS VDD _1925_ _1991_ _1992_ NOR2
X2873 VSS VDD _1925_ _1991_ _1892_ _1993_ OAI21
X2874 VSS VDD _1891_ _1993_ _1994_ NAND2
X2875 VSS VDD _1891_ _1993_ _1847_ _1995_ AOI21
X2876 VSS VDD _1846_ _1995_ _1996_ NOR2
X2877 VSS VDD _1695_ _1996_ _1684_ _1997_ OAI21
X2878 VSS VDD _1178_ _1200_ _1998_ XOR
X2879 VSS VDD _1998_ _1999_ INVERTER
X2880 VSS VDD _1997_ _1999_ _1211_ _2000_ AOI21
X2881 VSS VDD _0705_ _0804_ _2001_ XOR
X2882 VSS VDD _2000_ _2001_ _0815_ _2002_ OAI21
X2883 VSS VDD _0760_ _0793_ _2003_ NAND2
X2884 VSS VDD sensor4_6_ finestra_gaussiana4_6_ _0738_ _2004_ AOI21
X2885 VSS VDD _2003_ _2004_ _2005_ NAND2
X2886 VSS VDD _2003_ _2004_ _2006_ XOR
X2887 VSS VDD _2006_ _2007_ INVERTER
X2888 VSS VDD _2002_ _2006_ _2008_ NAND2
X2889 VSS VDD _0716_ _0727_ _2005_ _2008_ _2009_ OAI211
X2890 VSS VDD sensor5_7_ finestra_gaussiana5_3_ _2010_ NAND2
X2891 VSS VDD _2010_ _2011_ INVERTER
X2892 VSS VDD sensor5_6_ finestra_gaussiana5_4_ _2012_ NAND2
X2893 VSS VDD finestra_gaussiana5_5_ sensor5_5_ _2013_ NAND2
X2894 VSS VDD sensor5_6_ finestra_gaussiana5_5_ _2014_ NAND2
X2895 VSS VDD finestra_gaussiana5_4_ sensor5_5_ _2015_ NAND2
X2896 VSS VDD _2014_ _2015_ _2016_ NOR2
X2897 VSS VDD _2012_ _2013_ _2017_ XOR
X2898 VSS VDD _2011_ _2017_ _2018_ NAND2
X2899 VSS VDD sensor5_7_ finestra_gaussiana5_4_ _2019_ NAND2
X2900 VSS VDD sensor5_7_ finestra_gaussiana5_5_ _2020_ NAND2
X2901 VSS VDD _2012_ _2020_ _2021_ NOR2
X2902 VSS VDD _2014_ _2019_ _2022_ XOR
X2903 VSS VDD _2018_ _2022_ _2023_ XOR
X2904 VSS VDD finestra_gaussiana5_7_ sensor5_4_ _2024_ NAND2
X2905 VSS VDD finestra_gaussiana5_6_ _2016_ _2025_ NAND2
X2906 VSS VDD finestra_gaussiana5_6_ sensor5_5_ _2016_ _2026_ AOI21
X2907 VSS VDD finestra_gaussiana5_6_ _2016_ _2026_ _2027_ AOI21
X2908 VSS VDD finestra_gaussiana5_7_ sensor5_4_ _2027_ _2028_ AOI21
X2909 VSS VDD finestra_gaussiana5_6_ _2016_ _2024_ _2026_ _2029_ AOI211
X2910 VSS VDD finestra_gaussiana5_7_ sensor5_4_ _2027_ _2030_ NAND3
X2911 VSS VDD _2028_ _2029_ _2031_ NOR2
X2912 VSS VDD _2024_ _2027_ _2032_ XOR
X2913 VSS VDD _2023_ _2032_ _2033_ NOR2
X2914 VSS VDD _2011_ _2017_ _2022_ _2033_ _2034_ AOI31
X2915 VSS VDD finestra_gaussiana5_7_ sensor5_5_ _2035_ NAND2
X2916 VSS VDD finestra_gaussiana5_6_ _2021_ _2036_ NAND2
X2917 VSS VDD sensor5_6_ finestra_gaussiana5_6_ _2037_ NAND2
X2918 VSS VDD sensor5_6_ finestra_gaussiana5_6_ _2021_ _2038_ AOI21
X2919 VSS VDD _2012_ _2020_ _2037_ _2039_ OAI21
X2920 VSS VDD finestra_gaussiana5_6_ _2021_ _2038_ _2040_ AOI21
X2921 VSS VDD _2036_ _2039_ _2041_ NAND2
X2922 VSS VDD _2035_ _2041_ _2042_ XOR
X2923 VSS VDD _2035_ _2040_ _2043_ XOR
X2924 VSS VDD _2020_ _2043_ _2044_ NOR2
X2925 VSS VDD _2020_ _2043_ _2045_ XOR
X2926 VSS VDD _2020_ _2042_ _2046_ XOR
X2927 VSS VDD _2034_ _2046_ _2047_ NOR2
X2928 VSS VDD _2034_ _2045_ _2048_ XOR
X2929 VSS VDD _2024_ _2026_ _2025_ _2049_ OAI21
X2930 VSS VDD _2025_ _2030_ _2048_ _2050_ AOI21
X2931 VSS VDD _2047_ _2050_ _2051_ NOR2
X2932 VSS VDD finestra_gaussiana5_6_ sensor5_7_ _2052_ NAND2
X2933 VSS VDD finestra_gaussiana5_7_ sensor5_6_ _2053_ NAND2
X2934 VSS VDD finestra_gaussiana5_7_ sensor5_7_ _2054_ NAND2
X2935 VSS VDD _2052_ _2053_ _2055_ XOR
X2936 VSS VDD _2044_ _2055_ _2056_ NAND2
X2937 VSS VDD _2044_ _2055_ _2057_ XOR
X2938 VSS VDD _2035_ _2038_ _2036_ _2058_ OAI21
X2939 VSS VDD _2057_ _2058_ _2059_ NAND2
X2940 VSS VDD _2057_ _2058_ _2060_ XOR
X2941 VSS VDD _2047_ _2050_ _2060_ _2061_ OAI21
X2942 VSS VDD sensor5_5_ finestra_gaussiana5_3_ _2062_ NAND2
X2943 VSS VDD sensor5_7_ finestra_gaussiana5_1_ _2063_ NAND2
X2944 VSS VDD sensor5_5_ finestra_gaussiana5_1_ _2064_ NAND2
X2945 VSS VDD _2010_ _2064_ _2065_ NOR2
X2946 VSS VDD sensor5_6_ _2065_ _2066_ NAND2
X2947 VSS VDD sensor5_6_ finestra_gaussiana5_3_ _2067_ NAND2
X2948 VSS VDD _2010_ _2064_ _2067_ _2068_ OAI21
X2949 VSS VDD _2066_ _2068_ _2069_ NAND2
X2950 VSS VDD finestra_gaussiana5_5_ sensor5_4_ _2070_ NAND2
X2951 VSS VDD sensor5_7_ finestra_gaussiana5_2_ _2071_ NAND2
X2952 VSS VDD sensor5_5_ finestra_gaussiana5_2_ _2072_ NAND2
X2953 VSS VDD _2019_ _2072_ _2073_ NOR2
X2954 VSS VDD _2015_ _2071_ _2074_ XOR
X2955 VSS VDD _2070_ _2074_ _2075_ XOR
X2956 VSS VDD _2069_ _2075_ _2066_ _2076_ OAI21
X2957 VSS VDD _2011_ _2017_ _2077_ XOR
X2958 VSS VDD _2010_ _2017_ _2078_ XOR
X2959 VSS VDD _2076_ _2077_ _2079_ XOR
X2960 VSS VDD _2076_ _2078_ _2080_ XOR
X2961 VSS VDD finestra_gaussiana5_7_ sensor5_3_ _2081_ NAND2
X2962 VSS VDD finestra_gaussiana5_6_ sensor5_4_ _2082_ NAND2
X2963 VSS VDD finestra_gaussiana5_5_ sensor5_4_ _2074_ _2073_ _2083_ AOI31
X2964 VSS VDD _2082_ _2083_ _2084_ XOR
X2965 VSS VDD finestra_gaussiana5_7_ sensor5_3_ _2084_ _2085_ NAND3
X2966 VSS VDD _2081_ _2084_ _2086_ XOR
X2967 VSS VDD _2080_ _2086_ _2087_ NOR2
X2968 VSS VDD _2076_ _2077_ _2087_ _2088_ AOI21
X2969 VSS VDD _2023_ _2031_ _2089_ XOR
X2970 VSS VDD _2088_ _2089_ _2090_ NOR2
X2971 VSS VDD _2088_ _2089_ _2091_ XOR
X2972 VSS VDD _2082_ _2083_ _2085_ _2092_ OAI21
X2973 VSS VDD _2091_ _2092_ _2090_ _2093_ AOI21
X2974 VSS VDD _2048_ _2049_ _2094_ XOR
X2975 VSS VDD _2093_ _2094_ _2095_ NOR2
X2976 VSS VDD sensor5_7_ finestra_gaussiana5_0_ _2096_ NAND2
X2977 VSS VDD finestra_gaussiana5_3_ sensor5_4_ _2097_ NAND2
X2978 VSS VDD sensor5_4_ finestra_gaussiana5_0_ _2098_ NAND2
X2979 VSS VDD _2010_ _2098_ _2099_ NOR2
X2980 VSS VDD _2096_ _2097_ _2100_ XOR
X2981 VSS VDD sensor5_6_ finestra_gaussiana5_1_ _2101_ NAND2
X2982 VSS VDD sensor5_6_ finestra_gaussiana5_1_ _2100_ _2102_ NAND3
X2983 VSS VDD sensor5_6_ finestra_gaussiana5_1_ _2100_ _2099_ _2103_ AOI31
X2984 VSS VDD _2010_ _2098_ _2102_ _2104_ OAI21
X2985 VSS VDD _2062_ _2063_ _2105_ XOR
X2986 VSS VDD _2104_ _2105_ _2106_ NAND2
X2987 VSS VDD _2103_ _2105_ _2107_ XOR
X2988 VSS VDD finestra_gaussiana5_5_ sensor5_3_ _2108_ NAND2
X2989 VSS VDD finestra_gaussiana5_4_ sensor5_4_ _2109_ NAND2
X2990 VSS VDD sensor5_6_ finestra_gaussiana5_2_ _2110_ NAND2
X2991 VSS VDD sensor5_4_ finestra_gaussiana5_2_ _2111_ NAND2
X2992 VSS VDD _2012_ _2111_ _2112_ NOR2
X2993 VSS VDD _2109_ _2110_ _2113_ XOR
X2994 VSS VDD finestra_gaussiana5_5_ sensor5_3_ _2113_ _2114_ NAND3
X2995 VSS VDD _2108_ _2113_ _2115_ XOR
X2996 VSS VDD _2107_ _2115_ _2106_ _2116_ OAI21
X2997 VSS VDD _2069_ _2075_ _2117_ XOR
X2998 VSS VDD _2116_ _2117_ _2118_ NAND2
X2999 VSS VDD _2116_ _2117_ _2119_ XOR
X3000 VSS VDD finestra_gaussiana5_7_ sensor5_2_ _2120_ NAND2
X3001 VSS VDD finestra_gaussiana5_6_ sensor5_3_ _2121_ NAND2
X3002 VSS VDD finestra_gaussiana5_5_ sensor5_3_ _2113_ _2112_ _2122_ AOI31
X3003 VSS VDD _2012_ _2111_ _2114_ _2123_ OAI21
X3004 VSS VDD finestra_gaussiana5_6_ sensor5_3_ _2123_ _2124_ NAND3
X3005 VSS VDD _2121_ _2122_ _2125_ XOR
X3006 VSS VDD _2121_ _2123_ _2126_ XOR
X3007 VSS VDD finestra_gaussiana5_7_ sensor5_2_ _2125_ _2127_ NAND3
X3008 VSS VDD _2120_ _2126_ _2128_ XOR
X3009 VSS VDD _2120_ _2125_ _2129_ XOR
X3010 VSS VDD _2119_ _2128_ _2130_ NAND2
X3011 VSS VDD _2118_ _2130_ _2131_ NAND2
X3012 VSS VDD _2079_ _2086_ _2132_ XOR
X3013 VSS VDD _2118_ _2130_ _2132_ _2133_ AOI21
X3014 VSS VDD _2131_ _2132_ _2134_ XOR
X3015 VSS VDD _2124_ _2127_ _2135_ NAND2
X3016 VSS VDD _2124_ _2127_ _2134_ _2136_ AOI21
X3017 VSS VDD _2133_ _2136_ _2137_ NOR2
X3018 VSS VDD _2091_ _2092_ _2138_ XOR
X3019 VSS VDD _2133_ _2136_ _2138_ _2139_ OAI21
X3020 VSS VDD _2137_ _2138_ _2140_ XOR
X3021 VSS VDD _2140_ _2141_ INVERTER
X3022 VSS VDD sensor5_6_ finestra_gaussiana5_0_ _2142_ NAND2
X3023 VSS VDD finestra_gaussiana5_3_ sensor5_3_ _2143_ NAND2
X3024 VSS VDD sensor5_3_ finestra_gaussiana5_0_ _2144_ NAND2
X3025 VSS VDD _2067_ _2144_ _2145_ NOR2
X3026 VSS VDD _2142_ _2143_ _2146_ XOR
X3027 VSS VDD sensor5_5_ finestra_gaussiana5_1_ _2146_ _2145_ _2147_ AOI31
X3028 VSS VDD _2100_ _2101_ _2148_ XOR
X3029 VSS VDD _2147_ _2148_ _2149_ XOR
X3030 VSS VDD finestra_gaussiana5_5_ sensor5_2_ _2150_ NAND2
X3031 VSS VDD finestra_gaussiana5_4_ sensor5_3_ _2151_ NAND2
X3032 VSS VDD finestra_gaussiana5_2_ sensor5_3_ _2152_ NAND2
X3033 VSS VDD _2015_ _2152_ _2153_ NOR2
X3034 VSS VDD _2072_ _2151_ _2154_ NAND2
X3035 VSS VDD _2072_ _2151_ _2155_ XOR
X3036 VSS VDD _2015_ _2152_ _2154_ _2156_ OAI21
X3037 VSS VDD finestra_gaussiana5_5_ sensor5_2_ _2155_ _2157_ NAND3
X3038 VSS VDD _2150_ _2156_ _2158_ XOR
X3039 VSS VDD _2149_ _2158_ _2159_ NAND2
X3040 VSS VDD _2147_ _2148_ _2159_ _2160_ OAI21
X3041 VSS VDD _2107_ _2115_ _2161_ XOR
X3042 VSS VDD _2160_ _2161_ _2162_ NAND2
X3043 VSS VDD _2160_ _2161_ _2163_ XOR
X3044 VSS VDD finestra_gaussiana5_7_ sensor5_1_ _2164_ NAND2
X3045 VSS VDD finestra_gaussiana5_6_ sensor5_2_ _2165_ NAND2
X3046 VSS VDD finestra_gaussiana5_5_ sensor5_2_ _2154_ _2153_ _2166_ AOI31
X3047 VSS VDD _2015_ _2152_ _2157_ _2167_ OAI21
X3048 VSS VDD _2165_ _2166_ _2168_ XOR
X3049 VSS VDD _2165_ _2167_ _2169_ XOR
X3050 VSS VDD finestra_gaussiana5_7_ sensor5_1_ _2168_ _2170_ NAND3
X3051 VSS VDD _2164_ _2169_ _2171_ XOR
X3052 VSS VDD _2164_ _2168_ _2172_ XOR
X3053 VSS VDD _2163_ _2171_ _2173_ NAND2
X3054 VSS VDD _2162_ _2173_ _2174_ NAND2
X3055 VSS VDD _2119_ _2129_ _2175_ XOR
X3056 VSS VDD _2162_ _2173_ _2175_ _2176_ AOI21
X3057 VSS VDD _2162_ _2173_ _2175_ _2177_ NAND3
X3058 VSS VDD _2174_ _2175_ _2178_ XOR
X3059 VSS VDD _2165_ _2166_ _2170_ _2179_ OAI21
X3060 VSS VDD _2179_ _2180_ INVERTER
X3061 VSS VDD _2177_ _2179_ _2176_ _2181_ AOI21
X3062 VSS VDD _2134_ _2135_ _2182_ XOR
X3063 VSS VDD _2181_ _2182_ _2183_ NOR2
X3064 VSS VDD _2181_ _2182_ _2184_ XOR
X3065 VSS VDD sensor5_5_ finestra_gaussiana5_0_ _2185_ NAND2
X3066 VSS VDD finestra_gaussiana5_3_ sensor5_2_ _2186_ NAND2
X3067 VSS VDD finestra_gaussiana5_0_ sensor5_2_ _2187_ NAND2
X3068 VSS VDD _2062_ _2187_ _2188_ NOR2
X3069 VSS VDD sensor5_4_ finestra_gaussiana5_1_ _2189_ NAND2
X3070 VSS VDD _2189_ _2190_ INVERTER
X3071 VSS VDD _2185_ _2186_ _2191_ XOR
X3072 VSS VDD _2190_ _2191_ _2188_ _2192_ AOI21
X3073 VSS VDD _2064_ _2146_ _2193_ XOR
X3074 VSS VDD _2192_ _2193_ _2194_ NOR2
X3075 VSS VDD _2192_ _2193_ _2195_ XOR
X3076 VSS VDD finestra_gaussiana5_5_ sensor5_1_ _2196_ NAND2
X3077 VSS VDD finestra_gaussiana5_4_ sensor5_2_ _2197_ NAND2
X3078 VSS VDD _2197_ _2198_ INVERTER
X3079 VSS VDD finestra_gaussiana5_2_ sensor5_2_ _2199_ NAND2
X3080 VSS VDD _2111_ _2197_ _2200_ NOR2
X3081 VSS VDD _2111_ _2197_ _2201_ NAND2
X3082 VSS VDD _2111_ _2198_ _2202_ XOR
X3083 VSS VDD _2196_ _2202_ _2203_ XOR
X3084 VSS VDD _2195_ _2203_ _2194_ _2204_ AOI21
X3085 VSS VDD _2204_ _2205_ INVERTER
X3086 VSS VDD _2149_ _2158_ _2206_ XOR
X3087 VSS VDD _2205_ _2206_ _2207_ NAND2
X3088 VSS VDD _2204_ _2206_ _2208_ XOR
X3089 VSS VDD finestra_gaussiana5_7_ sensor5_0_ _2209_ NAND2
X3090 VSS VDD finestra_gaussiana5_6_ sensor5_1_ _2210_ NAND2
X3091 VSS VDD finestra_gaussiana5_5_ sensor5_1_ _2201_ _2200_ _2211_ AOI31
X3092 VSS VDD _2210_ _2211_ _2212_ NOR2
X3093 VSS VDD _2210_ _2211_ _2213_ XOR
X3094 VSS VDD _2209_ _2213_ _2214_ XOR
X3095 VSS VDD _2208_ _2214_ _2207_ _2215_ OAI21
X3096 VSS VDD _2215_ _2216_ INVERTER
X3097 VSS VDD _2163_ _2171_ _2217_ XOR
X3098 VSS VDD _2163_ _2172_ _2218_ XOR
X3099 VSS VDD _2216_ _2218_ _2219_ NOR2
X3100 VSS VDD _2215_ _2217_ _2220_ XOR
X3101 VSS VDD _2215_ _2218_ _2221_ XOR
X3102 VSS VDD finestra_gaussiana5_7_ sensor5_0_ _2213_ _2212_ _2222_ AOI31
X3103 VSS VDD _2221_ _2222_ _2223_ NOR2
X3104 VSS VDD _2219_ _2223_ _2224_ NOR2
X3105 VSS VDD _2178_ _2180_ _2225_ XOR
X3106 VSS VDD _2178_ _2179_ _2226_ XOR
X3107 VSS VDD _2219_ _2223_ _2225_ _2227_ OAI21
X3108 VSS VDD _2224_ _2226_ _2228_ XOR
X3109 VSS VDD _2224_ _2225_ _2229_ XOR
X3110 VSS VDD finestra_gaussiana5_3_ sensor5_1_ _2230_ NAND2
X3111 VSS VDD finestra_gaussiana5_0_ sensor5_1_ _2231_ NAND2
X3112 VSS VDD _2097_ _2231_ _2232_ NOR2
X3113 VSS VDD finestra_gaussiana5_1_ sensor5_3_ _2233_ NAND2
X3114 VSS VDD _2233_ _2234_ INVERTER
X3115 VSS VDD _2098_ _2230_ _2235_ XOR
X3116 VSS VDD _2234_ _2235_ _2232_ _2236_ AOI21
X3117 VSS VDD _2190_ _2191_ _2237_ XOR
X3118 VSS VDD _2189_ _2191_ _2238_ XOR
X3119 VSS VDD _2236_ _2238_ _2239_ NOR2
X3120 VSS VDD _2236_ _2238_ _2240_ XOR
X3121 VSS VDD _2236_ _2237_ _2241_ XOR
X3122 VSS VDD finestra_gaussiana5_5_ sensor5_0_ _2242_ NAND2
X3123 VSS VDD _2242_ _2243_ INVERTER
X3124 VSS VDD finestra_gaussiana5_4_ sensor5_1_ _2244_ NAND2
X3125 VSS VDD finestra_gaussiana5_2_ sensor5_1_ _2245_ NAND2
X3126 VSS VDD _2151_ _2245_ _2246_ NOR2
X3127 VSS VDD _2152_ _2244_ _2247_ XOR
X3128 VSS VDD _2243_ _2247_ _2248_ NAND2
X3129 VSS VDD _2243_ _2247_ _2249_ XOR
X3130 VSS VDD _2242_ _2247_ _2250_ XOR
X3131 VSS VDD _2241_ _2250_ _2251_ NOR2
X3132 VSS VDD _2240_ _2249_ _2239_ _2252_ AOI21
X3133 VSS VDD _2195_ _2203_ _2253_ XOR
X3134 VSS VDD _2239_ _2251_ _2253_ _2254_ OAI21
X3135 VSS VDD _2252_ _2253_ _2255_ XOR
X3136 VSS VDD finestra_gaussiana5_6_ sensor5_0_ _2256_ NAND2
X3137 VSS VDD _2243_ _2247_ _2246_ _2257_ AOI21
X3138 VSS VDD _2151_ _2245_ _2248_ _2258_ OAI21
X3139 VSS VDD _2256_ _2257_ _2259_ NOR2
X3140 VSS VDD _2256_ _2257_ _2260_ XOR
X3141 VSS VDD _2256_ _2258_ _2261_ XOR
X3142 VSS VDD _2255_ _2261_ _2254_ _2262_ OAI21
X3143 VSS VDD _2208_ _2214_ _2263_ XOR
X3144 VSS VDD _2262_ _2263_ _2264_ NAND2
X3145 VSS VDD _2262_ _2263_ _2265_ XOR
X3146 VSS VDD _2259_ _2265_ _2266_ NAND2
X3147 VSS VDD _2264_ _2266_ _2267_ NAND2
X3148 VSS VDD _2221_ _2222_ _2268_ XOR
X3149 VSS VDD _2220_ _2222_ _2269_ XOR
X3150 VSS VDD _2264_ _2266_ _2269_ _2270_ AOI21
X3151 VSS VDD _2234_ _2235_ _2271_ XOR
X3152 VSS VDD _2233_ _2235_ _2272_ XOR
X3153 VSS VDD finestra_gaussiana5_3_ sensor5_0_ _2273_ NAND2
X3154 VSS VDD finestra_gaussiana5_0_ sensor5_0_ _2274_ NAND2
X3155 VSS VDD _2143_ _2274_ _2275_ NOR2
X3156 VSS VDD finestra_gaussiana5_1_ sensor5_2_ _2276_ NAND2
X3157 VSS VDD _2144_ _2273_ _2276_ _2277_ AOI21
X3158 VSS VDD _2275_ _2277_ _2278_ NOR2
X3159 VSS VDD _2272_ _2278_ _2279_ NOR2
X3160 VSS VDD _2272_ _2278_ _2280_ XOR
X3161 VSS VDD _2271_ _2278_ _2281_ XOR
X3162 VSS VDD finestra_gaussiana5_4_ sensor5_0_ _2282_ NAND2
X3163 VSS VDD finestra_gaussiana5_2_ sensor5_0_ _2283_ NAND2
X3164 VSS VDD _2197_ _2283_ _2284_ NOR2
X3165 VSS VDD finestra_gaussiana5_2_ sensor5_0_ _2198_ _2285_ NAND3
X3166 VSS VDD _2199_ _2282_ _2286_ XOR
X3167 VSS VDD _2286_ _2287_ INVERTER
X3168 VSS VDD _2281_ _2287_ _2288_ NOR2
X3169 VSS VDD _2280_ _2286_ _2279_ _2289_ AOI21
X3170 VSS VDD _2240_ _2249_ _2290_ XOR
X3171 VSS VDD _2279_ _2288_ _2290_ _2291_ OAI21
X3172 VSS VDD _2289_ _2290_ _2292_ XOR
X3173 VSS VDD _2285_ _2292_ _2291_ _2293_ OAI21
X3174 VSS VDD _2293_ _2294_ INVERTER
X3175 VSS VDD _2255_ _2260_ _2295_ XOR
X3176 VSS VDD _2294_ _2295_ _2296_ NOR2
X3177 VSS VDD _2259_ _2265_ _2297_ XOR
X3178 VSS VDD _2296_ _2297_ _2298_ NAND2
X3179 VSS VDD _2144_ _2273_ _2299_ XOR
X3180 VSS VDD finestra_gaussiana5_1_ sensor5_1_ _2300_ NAND2
X3181 VSS VDD _2231_ _2276_ _2299_ _2301_ NOR3
X3182 VSS VDD finestra_gaussiana5_1_ sensor5_2_ _2231_ _2302_ NAND3
X3183 VSS VDD _2299_ _2302_ _2303_ XOR
X3184 VSS VDD _2245_ _2303_ _2304_ NOR2
X3185 VSS VDD _2301_ _2304_ _2305_ NOR2
X3186 VSS VDD _2280_ _2286_ _2306_ XOR
X3187 VSS VDD _2281_ _2286_ _2307_ XOR
X3188 VSS VDD _2301_ _2304_ _2306_ _2308_ OAI21
X3189 VSS VDD _2285_ _2292_ _2309_ XOR
X3190 VSS VDD _2284_ _2292_ _2310_ XOR
X3191 VSS VDD _2301_ _2304_ _2306_ _2309_ _2311_ OAI211
X3192 VSS VDD _2293_ _2295_ _2312_ XOR
X3193 VSS VDD _2311_ _2312_ _2313_ NOR2
X3194 VSS VDD finestra_gaussiana5_1_ sensor5_0_ _2314_ NAND2
X3195 VSS VDD _2274_ _2300_ _2315_ NOR2
X3196 VSS VDD _2187_ _2300_ _2316_ XOR
X3197 VSS VDD _2315_ _2316_ _2317_ NAND2
X3198 VSS VDD _2315_ _2316_ _2318_ NOR2
X3199 VSS VDD _2315_ _2316_ _2319_ XOR
X3200 VSS VDD _2283_ _2318_ _2317_ _2320_ OAI21
X3201 VSS VDD _2245_ _2303_ _2321_ XOR
X3202 VSS VDD _2320_ _2321_ _2322_ NAND2
X3203 VSS VDD _2305_ _2307_ _2323_ XOR
X3204 VSS VDD _2305_ _2306_ _2324_ XOR
X3205 VSS VDD _2322_ _2324_ _2325_ NOR2
X3206 VSS VDD _2309_ _2325_ _2326_ NAND2
X3207 VSS VDD _2326_ _2327_ INVERTER
X3208 VSS VDD _2311_ _2312_ _2328_ XOR
X3209 VSS VDD _2327_ _2328_ _2313_ _2329_ AOI21
X3210 VSS VDD _2296_ _2297_ _2330_ NOR2
X3211 VSS VDD _2296_ _2297_ _2331_ XOR
X3212 VSS VDD _2329_ _2330_ _2298_ _2332_ OAI21
X3213 VSS VDD _2267_ _2268_ _2333_ XOR
X3214 VSS VDD _2332_ _2333_ _2270_ _2334_ AOI21
X3215 VSS VDD _2229_ _2334_ _2227_ _2335_ OAI21
X3216 VSS VDD _2184_ _2335_ _2183_ _2336_ AOI21
X3217 VSS VDD _2140_ _2336_ _2139_ _2337_ OAI21
X3218 VSS VDD _2093_ _2094_ _2338_ XOR
X3219 VSS VDD _2337_ _2338_ _2095_ _2339_ AOI21
X3220 VSS VDD _2051_ _2060_ _2340_ XOR
X3221 VSS VDD _2340_ _2341_ INVERTER
X3222 VSS VDD _2339_ _2340_ _2061_ _2342_ OAI21
X3223 VSS VDD _2056_ _2059_ _2343_ NAND2
X3224 VSS VDD sensor5_6_ finestra_gaussiana5_6_ _2054_ _2344_ AOI21
X3225 VSS VDD finestra_gaussiana5_7_ sensor5_7_ _2037_ _2345_ NAND3
X3226 VSS VDD _2343_ _2344_ _2346_ XOR
X3227 VSS VDD _2343_ _2345_ _2347_ XOR
X3228 VSS VDD _2342_ _2346_ _2348_ XOR
X3229 VSS VDD _2342_ _2347_ _2349_ XOR
X3230 VSS VDD sensor6_7_ finestra_gaussiana6_3_ _2350_ NAND2
X3231 VSS VDD sensor6_6_ finestra_gaussiana6_4_ _2351_ NAND2
X3232 VSS VDD finestra_gaussiana6_5_ sensor6_5_ _2352_ NAND2
X3233 VSS VDD finestra_gaussiana6_5_ sensor6_6_ _2353_ NAND2
X3234 VSS VDD finestra_gaussiana6_4_ sensor6_5_ _2354_ NAND2
X3235 VSS VDD _2353_ _2354_ _2355_ NOR2
X3236 VSS VDD _2351_ _2352_ _2356_ NAND2
X3237 VSS VDD _2351_ _2352_ _2357_ XOR
X3238 VSS VDD _2353_ _2354_ _2356_ _2358_ OAI21
X3239 VSS VDD _2350_ _2358_ _2359_ NOR2
X3240 VSS VDD sensor6_7_ finestra_gaussiana6_4_ _2360_ NAND2
X3241 VSS VDD sensor6_7_ finestra_gaussiana6_5_ _2361_ NAND2
X3242 VSS VDD _2351_ _2361_ _2362_ NOR2
X3243 VSS VDD _2353_ _2360_ _2363_ XOR
X3244 VSS VDD _2359_ _2363_ _2364_ NAND2
X3245 VSS VDD _2359_ _2363_ _2365_ XOR
X3246 VSS VDD finestra_gaussiana6_7_ sensor6_4_ _2366_ NAND2
X3247 VSS VDD finestra_gaussiana6_6_ _2355_ _2367_ NAND2
X3248 VSS VDD finestra_gaussiana6_6_ sensor6_5_ _2355_ _2368_ AOI21
X3249 VSS VDD finestra_gaussiana6_6_ _2355_ _2368_ _2369_ AOI21
X3250 VSS VDD finestra_gaussiana6_7_ sensor6_4_ _2369_ _2370_ AOI21
X3251 VSS VDD finestra_gaussiana6_6_ _2355_ _2366_ _2368_ _2371_ AOI211
X3252 VSS VDD _2370_ _2371_ _2372_ NOR2
X3253 VSS VDD _2366_ _2369_ _2373_ XOR
X3254 VSS VDD _2365_ _2372_ _2374_ NAND2
X3255 VSS VDD finestra_gaussiana6_7_ sensor6_5_ _2375_ NAND2
X3256 VSS VDD finestra_gaussiana6_6_ _2362_ _2376_ NAND2
X3257 VSS VDD finestra_gaussiana6_6_ sensor6_6_ _2377_ NAND2
X3258 VSS VDD finestra_gaussiana6_6_ sensor6_6_ _2362_ _2378_ AOI21
X3259 VSS VDD _2351_ _2361_ _2377_ _2379_ OAI21
X3260 VSS VDD finestra_gaussiana6_6_ _2362_ _2378_ _2380_ AOI21
X3261 VSS VDD _2376_ _2379_ _2381_ NAND2
X3262 VSS VDD _2375_ _2381_ _2382_ XOR
X3263 VSS VDD _2375_ _2380_ _2383_ XOR
X3264 VSS VDD _2361_ _2383_ _2384_ NOR2
X3265 VSS VDD _2361_ _2382_ _2385_ XOR
X3266 VSS VDD _2364_ _2374_ _2385_ _2386_ AOI21
X3267 VSS VDD _2386_ _2387_ INVERTER
X3268 VSS VDD _2364_ _2374_ _2385_ _2388_ NAND3
X3269 VSS VDD _2387_ _2388_ _2389_ NAND2
X3270 VSS VDD _2366_ _2368_ _2367_ _2390_ OAI21
X3271 VSS VDD _2387_ _2388_ _2390_ _2391_ NAND3
X3272 VSS VDD _2388_ _2390_ _2386_ _2392_ AOI21
X3273 VSS VDD _2387_ _2391_ _2393_ NAND2
X3274 VSS VDD finestra_gaussiana6_6_ sensor6_7_ _2394_ NAND2
X3275 VSS VDD finestra_gaussiana6_7_ sensor6_6_ _2395_ NAND2
X3276 VSS VDD sensor6_7_ finestra_gaussiana6_7_ _2396_ NAND2
X3277 VSS VDD _2394_ _2395_ _2397_ XOR
X3278 VSS VDD _2384_ _2397_ _2398_ NAND2
X3279 VSS VDD _2384_ _2397_ _2399_ XOR
X3280 VSS VDD _2375_ _2378_ _2376_ _2400_ OAI21
X3281 VSS VDD _2399_ _2400_ _2401_ NAND2
X3282 VSS VDD _2399_ _2400_ _2402_ XOR
X3283 VSS VDD _2393_ _2402_ _2403_ NAND2
X3284 VSS VDD sensor6_5_ finestra_gaussiana6_3_ _2404_ NAND2
X3285 VSS VDD sensor6_7_ finestra_gaussiana6_1_ _2405_ NAND2
X3286 VSS VDD sensor6_5_ finestra_gaussiana6_1_ _2406_ NAND2
X3287 VSS VDD _2350_ _2406_ _2407_ NOR2
X3288 VSS VDD sensor6_6_ _2407_ _2408_ NAND2
X3289 VSS VDD sensor6_6_ finestra_gaussiana6_3_ _2409_ NAND2
X3290 VSS VDD _2350_ _2406_ _2409_ _2410_ OAI21
X3291 VSS VDD _2408_ _2410_ _2411_ NAND2
X3292 VSS VDD finestra_gaussiana6_5_ sensor6_4_ _2412_ NAND2
X3293 VSS VDD sensor6_7_ finestra_gaussiana6_2_ _2413_ NAND2
X3294 VSS VDD sensor6_5_ finestra_gaussiana6_2_ _2414_ NAND2
X3295 VSS VDD _2360_ _2414_ _2415_ NOR2
X3296 VSS VDD _2354_ _2413_ _2416_ XOR
X3297 VSS VDD _2412_ _2416_ _2417_ XOR
X3298 VSS VDD _2411_ _2417_ _2408_ _2418_ OAI21
X3299 VSS VDD _2350_ _2358_ _2419_ XOR
X3300 VSS VDD _2350_ _2357_ _2420_ XOR
X3301 VSS VDD _2418_ _2419_ _2421_ XOR
X3302 VSS VDD _2418_ _2420_ _2422_ XOR
X3303 VSS VDD finestra_gaussiana6_7_ sensor6_3_ _2423_ NAND2
X3304 VSS VDD finestra_gaussiana6_6_ sensor6_4_ _2424_ NAND2
X3305 VSS VDD finestra_gaussiana6_5_ sensor6_4_ _2416_ _2415_ _2425_ AOI31
X3306 VSS VDD _2424_ _2425_ _2426_ XOR
X3307 VSS VDD finestra_gaussiana6_7_ sensor6_3_ _2426_ _2427_ NAND3
X3308 VSS VDD _2423_ _2426_ _2428_ XOR
X3309 VSS VDD _2422_ _2428_ _2429_ NOR2
X3310 VSS VDD _2418_ _2419_ _2429_ _2430_ AOI21
X3311 VSS VDD _2365_ _2373_ _2431_ XOR
X3312 VSS VDD _2430_ _2431_ _2432_ NOR2
X3313 VSS VDD _2430_ _2431_ _2433_ XOR
X3314 VSS VDD _2424_ _2425_ _2427_ _2434_ OAI21
X3315 VSS VDD _2433_ _2434_ _2432_ _2435_ AOI21
X3316 VSS VDD _2389_ _2390_ _2436_ XOR
X3317 VSS VDD _2435_ _2436_ _2437_ NOR2
X3318 VSS VDD sensor6_7_ finestra_gaussiana6_0_ _2438_ NAND2
X3319 VSS VDD finestra_gaussiana6_3_ sensor6_4_ _2439_ NAND2
X3320 VSS VDD sensor6_4_ finestra_gaussiana6_0_ _2440_ NAND2
X3321 VSS VDD _2350_ _2440_ _2441_ NOR2
X3322 VSS VDD _2438_ _2439_ _2442_ XOR
X3323 VSS VDD sensor6_6_ finestra_gaussiana6_1_ _2443_ NAND2
X3324 VSS VDD sensor6_6_ finestra_gaussiana6_1_ _2442_ _2444_ NAND3
X3325 VSS VDD sensor6_6_ finestra_gaussiana6_1_ _2442_ _2441_ _2445_ AOI31
X3326 VSS VDD _2350_ _2440_ _2444_ _2446_ OAI21
X3327 VSS VDD _2404_ _2405_ _2447_ XOR
X3328 VSS VDD _2446_ _2447_ _2448_ NAND2
X3329 VSS VDD _2445_ _2447_ _2449_ XOR
X3330 VSS VDD finestra_gaussiana6_5_ sensor6_3_ _2450_ NAND2
X3331 VSS VDD finestra_gaussiana6_4_ sensor6_4_ _2451_ NAND2
X3332 VSS VDD sensor6_6_ finestra_gaussiana6_2_ _2452_ NAND2
X3333 VSS VDD sensor6_4_ finestra_gaussiana6_2_ _2453_ NAND2
X3334 VSS VDD _2351_ _2453_ _2454_ NOR2
X3335 VSS VDD _2451_ _2452_ _2455_ XOR
X3336 VSS VDD finestra_gaussiana6_5_ sensor6_3_ _2455_ _2456_ NAND3
X3337 VSS VDD _2450_ _2455_ _2457_ XOR
X3338 VSS VDD _2449_ _2457_ _2448_ _2458_ OAI21
X3339 VSS VDD _2411_ _2417_ _2459_ XOR
X3340 VSS VDD _2458_ _2459_ _2460_ NAND2
X3341 VSS VDD _2458_ _2459_ _2461_ XOR
X3342 VSS VDD finestra_gaussiana6_7_ sensor6_2_ _2462_ NAND2
X3343 VSS VDD finestra_gaussiana6_6_ sensor6_3_ _2463_ NAND2
X3344 VSS VDD finestra_gaussiana6_5_ sensor6_3_ _2455_ _2454_ _2464_ AOI31
X3345 VSS VDD _2351_ _2453_ _2456_ _2465_ OAI21
X3346 VSS VDD finestra_gaussiana6_6_ sensor6_3_ _2465_ _2466_ NAND3
X3347 VSS VDD _2463_ _2464_ _2467_ XOR
X3348 VSS VDD _2463_ _2465_ _2468_ XOR
X3349 VSS VDD finestra_gaussiana6_7_ sensor6_2_ _2467_ _2469_ NAND3
X3350 VSS VDD _2462_ _2468_ _2470_ XOR
X3351 VSS VDD _2461_ _2470_ _2471_ NAND2
X3352 VSS VDD _2460_ _2471_ _2472_ NAND2
X3353 VSS VDD _2421_ _2428_ _2473_ XOR
X3354 VSS VDD _2460_ _2471_ _2473_ _2474_ AOI21
X3355 VSS VDD _2472_ _2473_ _2475_ XOR
X3356 VSS VDD _2466_ _2469_ _2476_ NAND2
X3357 VSS VDD _2466_ _2469_ _2475_ _2477_ AOI21
X3358 VSS VDD _2474_ _2477_ _2478_ NOR2
X3359 VSS VDD _2433_ _2434_ _2479_ XOR
X3360 VSS VDD _2474_ _2477_ _2479_ _2480_ OAI21
X3361 VSS VDD _2478_ _2479_ _2481_ XOR
X3362 VSS VDD _2481_ _2482_ INVERTER
X3363 VSS VDD sensor6_6_ finestra_gaussiana6_0_ _2483_ NAND2
X3364 VSS VDD finestra_gaussiana6_3_ sensor6_3_ _2484_ NAND2
X3365 VSS VDD sensor6_3_ finestra_gaussiana6_0_ _2485_ NAND2
X3366 VSS VDD _2409_ _2485_ _2486_ NOR2
X3367 VSS VDD _2483_ _2484_ _2487_ XOR
X3368 VSS VDD sensor6_5_ finestra_gaussiana6_1_ _2487_ _2486_ _2488_ AOI31
X3369 VSS VDD _2442_ _2443_ _2489_ XOR
X3370 VSS VDD _2488_ _2489_ _2490_ XOR
X3371 VSS VDD finestra_gaussiana6_5_ sensor6_2_ _2491_ NAND2
X3372 VSS VDD finestra_gaussiana6_4_ sensor6_3_ _2492_ NAND2
X3373 VSS VDD finestra_gaussiana6_2_ sensor6_3_ _2493_ NAND2
X3374 VSS VDD _2414_ _2492_ _2494_ NAND2
X3375 VSS VDD _2414_ _2492_ _2495_ XOR
X3376 VSS VDD _2354_ _2493_ _2494_ _2496_ OAI21
X3377 VSS VDD finestra_gaussiana6_5_ sensor6_2_ _2495_ _2497_ NAND3
X3378 VSS VDD _2491_ _2496_ _2498_ XOR
X3379 VSS VDD _2491_ _2495_ _2499_ XOR
X3380 VSS VDD _2490_ _2498_ _2500_ NAND2
X3381 VSS VDD _2488_ _2489_ _2500_ _2501_ OAI21
X3382 VSS VDD _2449_ _2457_ _2502_ XOR
X3383 VSS VDD _2501_ _2502_ _2503_ NAND2
X3384 VSS VDD _2501_ _2502_ _2504_ XOR
X3385 VSS VDD finestra_gaussiana6_7_ sensor6_1_ _2505_ NAND2
X3386 VSS VDD finestra_gaussiana6_6_ sensor6_2_ _2506_ NAND2
X3387 VSS VDD _2354_ _2493_ _2497_ _2507_ OAI21
X3388 VSS VDD finestra_gaussiana6_6_ sensor6_2_ _2507_ _2508_ NAND3
X3389 VSS VDD _2506_ _2507_ _2509_ XOR
X3390 VSS VDD _2505_ _2509_ _2510_ XOR
X3391 VSS VDD _2504_ _2510_ _2511_ NAND2
X3392 VSS VDD _2503_ _2511_ _2512_ NAND2
X3393 VSS VDD _2461_ _2470_ _2513_ XOR
X3394 VSS VDD _2512_ _2513_ _2514_ NAND2
X3395 VSS VDD _2512_ _2513_ _2515_ XOR
X3396 VSS VDD _2505_ _2509_ _2508_ _2516_ OAI21
X3397 VSS VDD _2515_ _2516_ _2517_ NAND2
X3398 VSS VDD _2514_ _2517_ _2518_ NAND2
X3399 VSS VDD _2475_ _2476_ _2519_ XOR
X3400 VSS VDD _2519_ _2520_ INVERTER
X3401 VSS VDD _2514_ _2517_ _2519_ _2521_ AOI21
X3402 VSS VDD _2518_ _2520_ _2522_ XOR
X3403 VSS VDD sensor6_5_ finestra_gaussiana6_0_ _2523_ NAND2
X3404 VSS VDD finestra_gaussiana6_3_ sensor6_2_ _2524_ NAND2
X3405 VSS VDD finestra_gaussiana6_0_ sensor6_2_ _2525_ NAND2
X3406 VSS VDD _2404_ _2525_ _2526_ NOR2
X3407 VSS VDD sensor6_4_ finestra_gaussiana6_1_ _2527_ NAND2
X3408 VSS VDD _2527_ _2528_ INVERTER
X3409 VSS VDD _2523_ _2524_ _2529_ XOR
X3410 VSS VDD _2528_ _2529_ _2526_ _2530_ AOI21
X3411 VSS VDD _2406_ _2487_ _2531_ XOR
X3412 VSS VDD _2530_ _2531_ _2532_ NOR2
X3413 VSS VDD _2530_ _2531_ _2533_ XOR
X3414 VSS VDD finestra_gaussiana6_5_ sensor6_1_ _2534_ NAND2
X3415 VSS VDD finestra_gaussiana6_4_ sensor6_2_ _2535_ NAND2
X3416 VSS VDD finestra_gaussiana6_2_ sensor6_2_ _2536_ NAND2
X3417 VSS VDD _2453_ _2535_ _2537_ XOR
X3418 VSS VDD finestra_gaussiana6_5_ sensor6_1_ _2537_ _2538_ NAND3
X3419 VSS VDD _2534_ _2537_ _2539_ XOR
X3420 VSS VDD _2539_ _2540_ INVERTER
X3421 VSS VDD _2533_ _2540_ _2532_ _2541_ AOI21
X3422 VSS VDD _2490_ _2499_ _2542_ XOR
X3423 VSS VDD _2541_ _2542_ _2543_ NOR2
X3424 VSS VDD _2541_ _2542_ _2544_ XOR
X3425 VSS VDD finestra_gaussiana6_7_ sensor6_0_ _2545_ NAND2
X3426 VSS VDD finestra_gaussiana6_6_ sensor6_1_ _2546_ NAND2
X3427 VSS VDD _2451_ _2536_ _2538_ _2547_ OAI21
X3428 VSS VDD _2546_ _2547_ _2548_ XOR
X3429 VSS VDD _2545_ _2548_ _2549_ NOR2
X3430 VSS VDD _2545_ _2548_ _2550_ XOR
X3431 VSS VDD _2544_ _2550_ _2551_ NAND2
X3432 VSS VDD _2544_ _2550_ _2543_ _2552_ AOI21
X3433 VSS VDD _2541_ _2542_ _2551_ _2553_ OAI21
X3434 VSS VDD _2504_ _2510_ _2554_ XOR
X3435 VSS VDD _2553_ _2554_ _2555_ NAND2
X3436 VSS VDD _2553_ _2554_ _0017_ XOR
X3437 VSS VDD _2552_ _2554_ _0018_ XOR
X3438 VSS VDD finestra_gaussiana6_6_ sensor6_1_ _2547_ _2549_ _0019_ AOI31
X3439 VSS VDD _0018_ _0019_ _0020_ NOR2
X3440 VSS VDD _2553_ _2554_ _0020_ _0021_ AOI21
X3441 VSS VDD _0018_ _0019_ _2555_ _0022_ OAI21
X3442 VSS VDD _2515_ _2516_ _0023_ XOR
X3443 VSS VDD _0022_ _0023_ _0024_ NAND2
X3444 VSS VDD _0022_ _0023_ _0025_ XOR
X3445 VSS VDD _0021_ _0023_ _0026_ XOR
X3446 VSS VDD finestra_gaussiana6_3_ sensor6_1_ _0027_ NAND2
X3447 VSS VDD finestra_gaussiana6_0_ sensor6_1_ _0028_ NAND2
X3448 VSS VDD _2439_ _0028_ _0029_ NOR2
X3449 VSS VDD finestra_gaussiana6_1_ sensor6_3_ _0030_ NAND2
X3450 VSS VDD _0030_ _0031_ INVERTER
X3451 VSS VDD _2440_ _0027_ _0032_ XOR
X3452 VSS VDD _0031_ _0032_ _0029_ _0033_ AOI21
X3453 VSS VDD _2528_ _2529_ _0034_ XOR
X3454 VSS VDD _2527_ _2529_ _0035_ XOR
X3455 VSS VDD _0033_ _0035_ _0036_ NOR2
X3456 VSS VDD _0033_ _0035_ _0037_ XOR
X3457 VSS VDD _0033_ _0034_ _0038_ XOR
X3458 VSS VDD finestra_gaussiana6_5_ sensor6_0_ _0039_ NAND2
X3459 VSS VDD _0039_ _0040_ INVERTER
X3460 VSS VDD finestra_gaussiana6_4_ sensor6_1_ _0041_ NAND2
X3461 VSS VDD finestra_gaussiana6_2_ sensor6_1_ _0042_ NAND2
X3462 VSS VDD _2492_ _0042_ _0043_ NOR2
X3463 VSS VDD _2493_ _0041_ _0044_ XOR
X3464 VSS VDD _0040_ _0044_ _0045_ NAND2
X3465 VSS VDD _0040_ _0044_ _0046_ XOR
X3466 VSS VDD _0039_ _0044_ _0047_ XOR
X3467 VSS VDD _0038_ _0047_ _0048_ NOR2
X3468 VSS VDD _0037_ _0046_ _0036_ _0049_ AOI21
X3469 VSS VDD _2533_ _2540_ _0050_ XOR
X3470 VSS VDD _0036_ _0048_ _0050_ _0051_ OAI21
X3471 VSS VDD _0049_ _0050_ _0052_ XOR
X3472 VSS VDD finestra_gaussiana6_6_ sensor6_0_ _0053_ NAND2
X3473 VSS VDD _0040_ _0044_ _0043_ _0054_ AOI21
X3474 VSS VDD _2492_ _0042_ _0045_ _0055_ OAI21
X3475 VSS VDD _0053_ _0054_ _0056_ NOR2
X3476 VSS VDD _0053_ _0054_ _0057_ XOR
X3477 VSS VDD _0053_ _0055_ _0058_ XOR
X3478 VSS VDD _0052_ _0058_ _0051_ _0059_ OAI21
X3479 VSS VDD _2544_ _2550_ _0060_ XOR
X3480 VSS VDD _0059_ _0060_ _0061_ NAND2
X3481 VSS VDD _0059_ _0060_ _0062_ XOR
X3482 VSS VDD _0056_ _0062_ _0063_ NAND2
X3483 VSS VDD _0061_ _0063_ _0064_ NAND2
X3484 VSS VDD _0018_ _0019_ _0065_ XOR
X3485 VSS VDD _0017_ _0019_ _0066_ XOR
X3486 VSS VDD _0061_ _0063_ _0066_ _0067_ AOI21
X3487 VSS VDD _0031_ _0032_ _0068_ XOR
X3488 VSS VDD _0030_ _0032_ _0069_ XOR
X3489 VSS VDD finestra_gaussiana6_3_ sensor6_0_ _0070_ NAND2
X3490 VSS VDD finestra_gaussiana6_0_ sensor6_0_ _0071_ NAND2
X3491 VSS VDD _2484_ _0071_ _0072_ NOR2
X3492 VSS VDD finestra_gaussiana6_1_ sensor6_2_ _0073_ NAND2
X3493 VSS VDD _2485_ _0070_ _0073_ _0074_ AOI21
X3494 VSS VDD _0072_ _0074_ _0075_ NOR2
X3495 VSS VDD _0069_ _0075_ _0076_ NOR2
X3496 VSS VDD _0069_ _0075_ _0077_ XOR
X3497 VSS VDD _0068_ _0075_ _0078_ XOR
X3498 VSS VDD finestra_gaussiana6_4_ sensor6_0_ _0079_ NAND2
X3499 VSS VDD finestra_gaussiana6_2_ sensor6_0_ _0080_ NAND2
X3500 VSS VDD _0080_ _0081_ INVERTER
X3501 VSS VDD _2535_ _0080_ _0082_ NOR2
X3502 VSS VDD _2536_ _0079_ _0083_ XOR
X3503 VSS VDD _0083_ _0084_ INVERTER
X3504 VSS VDD _0078_ _0084_ _0085_ NOR2
X3505 VSS VDD _0077_ _0083_ _0076_ _0086_ AOI21
X3506 VSS VDD _0037_ _0046_ _0087_ XOR
X3507 VSS VDD _0076_ _0085_ _0087_ _0088_ OAI21
X3508 VSS VDD _0086_ _0087_ _0089_ XOR
X3509 VSS VDD _2535_ _0080_ _0088_ _0089_ _0090_ OAI31
X3510 VSS VDD _0090_ _0091_ INVERTER
X3511 VSS VDD _0052_ _0058_ _0092_ XOR
X3512 VSS VDD _0052_ _0057_ _0093_ XOR
X3513 VSS VDD _0091_ _0093_ _0094_ NOR2
X3514 VSS VDD _0090_ _0092_ _0095_ NAND2
X3515 VSS VDD _0056_ _0062_ _0096_ XOR
X3516 VSS VDD _0094_ _0096_ _0097_ NAND2
X3517 VSS VDD _0094_ _0096_ _0098_ XOR
X3518 VSS VDD _0095_ _0096_ _0099_ XOR
X3519 VSS VDD _2485_ _0070_ _0100_ XOR
X3520 VSS VDD finestra_gaussiana6_1_ sensor6_1_ _0101_ NAND2
X3521 VSS VDD finestra_gaussiana6_0_ sensor6_1_ _0073_ _0102_ AOI21
X3522 VSS VDD finestra_gaussiana6_1_ sensor6_2_ _0028_ _0103_ NAND3
X3523 VSS VDD _0100_ _0103_ _0104_ XOR
X3524 VSS VDD _0100_ _0102_ _0105_ XOR
X3525 VSS VDD finestra_gaussiana6_2_ sensor6_1_ _0105_ _0106_ NAND3
X3526 VSS VDD _0028_ _0073_ _0106_ _0100_ _0107_ OAI31
X3527 VSS VDD _0077_ _0083_ _0108_ XOR
X3528 VSS VDD _0078_ _0083_ _0109_ XOR
X3529 VSS VDD _0107_ _0108_ _0110_ NAND2
X3530 VSS VDD _0082_ _0089_ _0111_ XOR
X3531 VSS VDD _0110_ _0111_ _0112_ NOR2
X3532 VSS VDD _0090_ _0093_ _0113_ XOR
X3533 VSS VDD _0110_ _0111_ _0113_ _0114_ NOR3
X3534 VSS VDD finestra_gaussiana6_1_ sensor6_0_ _0115_ NAND2
X3535 VSS VDD _0071_ _0101_ _0116_ NOR2
X3536 VSS VDD _2525_ _0101_ _0117_ XOR
X3537 VSS VDD _0116_ _0117_ _0118_ NAND2
X3538 VSS VDD _0116_ _0117_ _0119_ NOR2
X3539 VSS VDD _0116_ _0117_ _0120_ XOR
X3540 VSS VDD _0080_ _0119_ _0118_ _0121_ OAI21
X3541 VSS VDD _0042_ _0104_ _0122_ XOR
X3542 VSS VDD _0121_ _0122_ _0123_ NAND2
X3543 VSS VDD _0107_ _0108_ _0124_ XOR
X3544 VSS VDD _0107_ _0109_ _0125_ XOR
X3545 VSS VDD _0123_ _0125_ _0126_ NOR2
X3546 VSS VDD _0121_ _0122_ _0124_ _0127_ NAND3
X3547 VSS VDD _0110_ _0111_ _0128_ XOR
X3548 VSS VDD _0126_ _0128_ _0129_ NAND2
X3549 VSS VDD _0110_ _0111_ _0113_ _0130_ OAI21
X3550 VSS VDD _0112_ _0113_ _0131_ XOR
X3551 VSS VDD _0126_ _0128_ _0130_ _0114_ _0132_ AOI31
X3552 VSS VDD _0099_ _0132_ _0097_ _0133_ OAI21
X3553 VSS VDD _0064_ _0065_ _0134_ XOR
X3554 VSS VDD _0064_ _0066_ _0135_ XOR
X3555 VSS VDD _0133_ _0134_ _0067_ _0136_ AOI21
X3556 VSS VDD _0026_ _0136_ _0024_ _0137_ OAI21
X3557 VSS VDD _2522_ _0137_ _2521_ _0138_ AOI21
X3558 VSS VDD _2481_ _0138_ _2480_ _0139_ OAI21
X3559 VSS VDD _2435_ _2436_ _0140_ XOR
X3560 VSS VDD _0139_ _0140_ _2437_ _0141_ AOI21
X3561 VSS VDD _2393_ _2402_ _0142_ XOR
X3562 VSS VDD _2392_ _2402_ _0143_ XOR
X3563 VSS VDD _0141_ _0143_ _2403_ _0144_ OAI21
X3564 VSS VDD _2398_ _2401_ _0145_ NAND2
X3565 VSS VDD finestra_gaussiana6_6_ sensor6_6_ _2396_ _0146_ AOI21
X3566 VSS VDD _0145_ _0146_ _0147_ XOR
X3567 VSS VDD _0144_ _0147_ _0148_ XOR
X3568 VSS VDD _2348_ _0148_ _0149_ NAND2
X3569 VSS VDD _2339_ _2341_ _0150_ XOR
X3570 VSS VDD _0141_ _0143_ _0151_ XOR
X3571 VSS VDD _0141_ _0142_ _0152_ XOR
X3572 VSS VDD _0150_ _0152_ _0153_ NOR2
X3573 VSS VDD _2337_ _2338_ _0154_ XOR
X3574 VSS VDD _0139_ _0140_ _0155_ XOR
X3575 VSS VDD _0154_ _0155_ _0156_ NAND2
X3576 VSS VDD _2141_ _2336_ _0157_ XOR
X3577 VSS VDD _2481_ _0138_ _0158_ XOR
X3578 VSS VDD _2482_ _0138_ _0159_ XOR
X3579 VSS VDD _0157_ _0159_ _0160_ NOR2
X3580 VSS VDD _0157_ _0159_ _0161_ XOR
X3581 VSS VDD _0157_ _0158_ _0162_ XOR
X3582 VSS VDD _2184_ _2335_ _0163_ XOR
X3583 VSS VDD _2522_ _0137_ _0164_ XOR
X3584 VSS VDD _0163_ _0164_ _0165_ NAND2
X3585 VSS VDD _2228_ _2334_ _0166_ XOR
X3586 VSS VDD _0026_ _0136_ _0167_ XOR
X3587 VSS VDD _0025_ _0136_ _0168_ XOR
X3588 VSS VDD _0166_ _0168_ _0169_ NOR2
X3589 VSS VDD _0166_ _0168_ _0170_ XOR
X3590 VSS VDD _0166_ _0167_ _0171_ XOR
X3591 VSS VDD _2332_ _2333_ _0172_ XOR
X3592 VSS VDD _0133_ _0134_ _0173_ XOR
X3593 VSS VDD _0133_ _0135_ _0174_ XOR
X3594 VSS VDD _0172_ _0173_ _0175_ NAND2
X3595 VSS VDD _2329_ _2331_ _0176_ XOR
X3596 VSS VDD _0099_ _0132_ _0177_ XOR
X3597 VSS VDD _0098_ _0132_ _0178_ XOR
X3598 VSS VDD _0176_ _0178_ _0179_ NOR2
X3599 VSS VDD _0176_ _0178_ _0180_ XOR
X3600 VSS VDD _0176_ _0177_ _0181_ XOR
X3601 VSS VDD _2327_ _2328_ _0182_ XOR
X3602 VSS VDD _2326_ _2328_ _0183_ XOR
X3603 VSS VDD _0129_ _0131_ _0184_ XOR
X3604 VSS VDD _0182_ _0184_ _0185_ NAND2
X3605 VSS VDD _0183_ _0184_ _0186_ XOR
X3606 VSS VDD _2322_ _2324_ _2308_ _0187_ OAI21
X3607 VSS VDD _2310_ _0187_ _0188_ XOR
X3608 VSS VDD _0127_ _0128_ _0189_ XOR
X3609 VSS VDD _0188_ _0189_ _0190_ NOR2
X3610 VSS VDD _0188_ _0189_ _0191_ XOR
X3611 VSS VDD _2322_ _2323_ _0192_ XOR
X3612 VSS VDD _0123_ _0124_ _0193_ XOR
X3613 VSS VDD _0192_ _0193_ _0194_ NOR2
X3614 VSS VDD _2320_ _2321_ _0195_ XOR
X3615 VSS VDD _0121_ _0122_ _0196_ XOR
X3616 VSS VDD _0195_ _0196_ _0197_ NAND2
X3617 VSS VDD _2283_ _2319_ _0198_ XOR
X3618 VSS VDD _0081_ _0120_ _0199_ XOR
X3619 VSS VDD _0080_ _0120_ _0200_ XOR
X3620 VSS VDD _0198_ _0200_ _0201_ NOR2
X3621 VSS VDD _2231_ _2314_ _0202_ XOR
X3622 VSS VDD _0028_ _0115_ _0203_ XOR
X3623 VSS VDD _0202_ _0203_ _0204_ NAND2
X3624 VSS VDD _2274_ _0071_ _0205_ NOR2
X3625 VSS VDD _0202_ _0203_ _0206_ NOR2
X3626 VSS VDD _0202_ _0203_ _0207_ XOR
X3627 VSS VDD _2274_ _0071_ _0204_ _0206_ _0208_ OAI31
X3628 VSS VDD _0198_ _0200_ _0209_ XOR
X3629 VSS VDD _0198_ _0199_ _0210_ XOR
X3630 VSS VDD _0208_ _0209_ _0201_ _0211_ AOI21
X3631 VSS VDD _0195_ _0196_ _0212_ NOR2
X3632 VSS VDD _0195_ _0196_ _0213_ XOR
X3633 VSS VDD _0211_ _0212_ _0197_ _0214_ OAI21
X3634 VSS VDD _0192_ _0193_ _0215_ XOR
X3635 VSS VDD _0214_ _0215_ _0194_ _0216_ AOI21
X3636 VSS VDD _0216_ _0217_ INVERTER
X3637 VSS VDD _0191_ _0217_ _0190_ _0218_ AOI21
X3638 VSS VDD _0186_ _0218_ _0185_ _0219_ OAI21
X3639 VSS VDD _0180_ _0219_ _0179_ _0220_ AOI21
X3640 VSS VDD _0172_ _0174_ _0221_ XOR
X3641 VSS VDD _0220_ _0221_ _0175_ _0222_ OAI21
X3642 VSS VDD _0170_ _0222_ _0169_ _0223_ AOI21
X3643 VSS VDD _0163_ _0164_ _0224_ NOR2
X3644 VSS VDD _0163_ _0164_ _0225_ XOR
X3645 VSS VDD _0223_ _0224_ _0165_ _0226_ OAI21
X3646 VSS VDD _0161_ _0226_ _0160_ _0227_ AOI21
X3647 VSS VDD _0154_ _0155_ _0228_ NOR2
X3648 VSS VDD _0154_ _0155_ _0229_ XOR
X3649 VSS VDD _0227_ _0228_ _0156_ _0230_ OAI21
X3650 VSS VDD _0150_ _0152_ _0231_ XOR
X3651 VSS VDD _0150_ _0151_ _0232_ XOR
X3652 VSS VDD _0230_ _0231_ _0153_ _0233_ AOI21
X3653 VSS VDD _2348_ _0148_ _0234_ XOR
X3654 VSS VDD _2349_ _0148_ _0235_ XOR
X3655 VSS VDD _0233_ _0235_ _0149_ _0236_ OAI21
X3656 VSS VDD _2037_ _2056_ _2059_ _2054_ _0237_ AOI31
X3657 VSS VDD _2342_ _2346_ _0237_ _0238_ AOI21
X3658 VSS VDD _2377_ _2398_ _2401_ _2396_ _0239_ AOI31
X3659 VSS VDD _0144_ _0147_ _0239_ _0240_ AOI21
X3660 VSS VDD _0238_ _0240_ _0241_ NOR2
X3661 VSS VDD _0238_ _0240_ _0242_ XOR
X3662 VSS VDD _0236_ _0242_ _0243_ XOR
X3663 VSS VDD _2002_ _2007_ _0244_ XOR
X3664 VSS VDD _0233_ _0235_ _0245_ XOR
X3665 VSS VDD _0233_ _0234_ _0246_ XOR
X3666 VSS VDD _0244_ _0246_ _0247_ NOR2
X3667 VSS VDD _2000_ _2001_ _0248_ XOR
X3668 VSS VDD _0230_ _0231_ _0249_ XOR
X3669 VSS VDD _0230_ _0232_ _0250_ XOR
X3670 VSS VDD _0248_ _0249_ _0251_ NAND2
X3671 VSS VDD _0248_ _0250_ _0252_ XOR
X3672 VSS VDD _1997_ _1999_ _0253_ XOR
X3673 VSS VDD _1997_ _1998_ _0254_ XOR
X3674 VSS VDD _0227_ _0229_ _0255_ XOR
X3675 VSS VDD _0254_ _0255_ _0256_ NOR2
X3676 VSS VDD _0254_ _0255_ _0257_ XOR
X3677 VSS VDD _0253_ _0255_ _0258_ XOR
X3678 VSS VDD _1695_ _1996_ _0259_ XOR
X3679 VSS VDD _0161_ _0226_ _0260_ XOR
X3680 VSS VDD _0162_ _0226_ _0261_ XOR
X3681 VSS VDD _0259_ _0260_ _0262_ NOR2
X3682 VSS VDD _0259_ _0260_ _0263_ NAND2
X3683 VSS VDD _1847_ _1994_ _0264_ XOR
X3684 VSS VDD _0223_ _0225_ _0265_ XOR
X3685 VSS VDD _0264_ _0265_ _0266_ NOR2
X3686 VSS VDD _0264_ _0265_ _0267_ XOR
X3687 VSS VDD _1893_ _1992_ _0268_ XOR
X3688 VSS VDD _1892_ _1992_ _0269_ XOR
X3689 VSS VDD _0170_ _0222_ _0270_ XOR
X3690 VSS VDD _0171_ _0222_ _0271_ XOR
X3691 VSS VDD _0269_ _0271_ _0272_ NOR2
X3692 VSS VDD _0268_ _0270_ _0273_ NAND2
X3693 VSS VDD _0269_ _0271_ _0274_ NAND2
X3694 VSS VDD _1988_ _1990_ _0275_ XOR
X3695 VSS VDD _1988_ _1989_ _0276_ XOR
X3696 VSS VDD _0220_ _0221_ _0277_ XOR
X3697 VSS VDD _0275_ _0277_ _0278_ NAND2
X3698 VSS VDD _1984_ _1986_ _0279_ XOR
X3699 VSS VDD _0181_ _0219_ _0280_ XOR
X3700 VSS VDD _0279_ _0280_ _0281_ NOR2
X3701 VSS VDD _0279_ _0280_ _0282_ XOR
X3702 VSS VDD _1982_ _1983_ _0283_ XOR
X3703 VSS VDD _0186_ _0218_ _0284_ XOR
X3704 VSS VDD _0283_ _0284_ _0285_ NAND2
X3705 VSS VDD _0283_ _0284_ _0286_ NOR2
X3706 VSS VDD _0283_ _0284_ _0288_ XOR
X3707 VSS VDD _0191_ _0216_ _0289_ XOR
X3708 VSS VDD _1979_ _1980_ _1963_ _0290_ OAI21
X3709 VSS VDD _1964_ _0290_ _0291_ XOR
X3710 VSS VDD _1965_ _0290_ _0292_ XOR
X3711 VSS VDD _0289_ _0292_ _0293_ NOR2
X3712 VSS VDD _0289_ _0292_ _0294_ NAND2
X3713 VSS VDD _0289_ _0291_ _0295_ XOR
X3714 VSS VDD _1979_ _1980_ _0296_ XOR
X3715 VSS VDD _0214_ _0215_ _0297_ XOR
X3716 VSS VDD _0296_ _0297_ _0299_ NAND2
X3717 VSS VDD _1976_ _1978_ _0300_ XOR
X3718 VSS VDD _0211_ _0213_ _0301_ XOR
X3719 VSS VDD _0300_ _0301_ _0302_ NOR2
X3720 VSS VDD _0300_ _0301_ _0303_ XOR
X3721 VSS VDD _1935_ _1975_ _0304_ XOR
X3722 VSS VDD _0208_ _0209_ _0305_ XOR
X3723 VSS VDD _0208_ _0210_ _0306_ XOR
X3724 VSS VDD _0304_ _0306_ _0307_ NOR2
X3725 VSS VDD _1895_ _1970_ _0308_ XOR
X3726 VSS VDD _0205_ _0207_ _0310_ XOR
X3727 VSS VDD _0308_ _0310_ _0311_ NAND2
X3728 VSS VDD _2274_ _0071_ _0312_ XOR
X3729 VSS VDD _0312_ _0313_ INVERTER
X3730 VSS VDD _1928_ _0313_ _0314_ NOR2
X3731 VSS VDD _0308_ _0310_ _0315_ NOR2
X3732 VSS VDD _0308_ _0310_ _0316_ XOR
X3733 VSS VDD _1928_ _0315_ _0311_ _0313_ _0317_ OAI31
X3734 VSS VDD _0304_ _0306_ _0318_ XOR
X3735 VSS VDD _0304_ _0305_ _0319_ XOR
X3736 VSS VDD _0317_ _0318_ _0321_ NAND2
X3737 VSS VDD _0317_ _0318_ _0307_ _0322_ AOI21
X3738 VSS VDD _0304_ _0306_ _0321_ _0323_ OAI21
X3739 VSS VDD _0303_ _0323_ _0302_ _0324_ AOI21
X3740 VSS VDD _0296_ _0297_ _0325_ NOR2
X3741 VSS VDD _0296_ _0297_ _0326_ XOR
X3742 VSS VDD _0324_ _0325_ _0299_ _0327_ OAI21
X3743 VSS VDD _0327_ _0328_ INVERTER
X3744 VSS VDD _0294_ _0327_ _0293_ _0329_ AOI21
X3745 VSS VDD _0286_ _0329_ _0285_ _0330_ OAI21
X3746 VSS VDD _0282_ _0330_ _0281_ _0332_ AOI21
X3747 VSS VDD _0275_ _0277_ _0333_ XOR
X3748 VSS VDD _0276_ _0277_ _0334_ XOR
X3749 VSS VDD _0332_ _0334_ _0278_ _0335_ OAI21
X3750 VSS VDD _0332_ _0334_ _0273_ _0278_ _0336_ OAI211
X3751 VSS VDD _0272_ _0335_ _0274_ _0337_ OAI21
X3752 VSS VDD _0267_ _0274_ _0336_ _0266_ _0338_ AOI31
X3753 VSS VDD _0262_ _0338_ _0263_ _0339_ OAI21
X3754 VSS VDD _0257_ _0339_ _0256_ _0340_ AOI21
X3755 VSS VDD _0252_ _0340_ _0251_ _0341_ OAI21
X3756 VSS VDD _0244_ _0246_ _0343_ XOR
X3757 VSS VDD _0244_ _0245_ _0344_ XOR
X3758 VSS VDD _0341_ _0343_ _0247_ _0345_ AOI21
X3759 VSS VDD _2009_ _0243_ _0346_ XOR
X3760 VSS VDD _0346_ _0347_ INVERTER
X3761 VSS VDD _0345_ _0347_ _0348_ NOR2
X3762 VSS VDD _2009_ _0243_ _0348_ _0349_ AOI21
X3763 VSS VDD _0236_ _0242_ _0241_ _0350_ AOI21
X3764 VSS VDD _0350_ _0351_ INVERTER
X3765 VSS VDD _0349_ _0350_ _0352_ NOR2
X3766 VSS VDD sensor2_7_ finestra_gaussiana2_3_ _0354_ NAND2
X3767 VSS VDD _0354_ _0355_ INVERTER
X3768 VSS VDD sensor2_6_ finestra_gaussiana2_4_ _0356_ NAND2
X3769 VSS VDD finestra_gaussiana2_5_ sensor2_5_ _0357_ NAND2
X3770 VSS VDD sensor2_6_ finestra_gaussiana2_5_ _0358_ NAND2
X3771 VSS VDD finestra_gaussiana2_4_ sensor2_5_ _0359_ NAND2
X3772 VSS VDD _0358_ _0359_ _0360_ NOR2
X3773 VSS VDD _0356_ _0357_ _0361_ XOR
X3774 VSS VDD _0355_ _0361_ _0362_ NAND2
X3775 VSS VDD sensor2_7_ finestra_gaussiana2_4_ _0363_ NAND2
X3776 VSS VDD sensor2_7_ finestra_gaussiana2_5_ _0365_ NAND2
X3777 VSS VDD _0356_ _0365_ _0366_ NOR2
X3778 VSS VDD _0358_ _0363_ _0367_ XOR
X3779 VSS VDD _0362_ _0367_ _0368_ XOR
X3780 VSS VDD finestra_gaussiana2_7_ sensor2_4_ _0369_ NAND2
X3781 VSS VDD finestra_gaussiana2_6_ _0360_ _0370_ NAND2
X3782 VSS VDD finestra_gaussiana2_6_ sensor2_5_ _0360_ _0371_ AOI21
X3783 VSS VDD finestra_gaussiana2_6_ _0360_ _0371_ _0372_ AOI21
X3784 VSS VDD finestra_gaussiana2_7_ sensor2_4_ _0372_ _0373_ AOI21
X3785 VSS VDD finestra_gaussiana2_6_ _0360_ _0369_ _0371_ _0374_ AOI211
X3786 VSS VDD finestra_gaussiana2_7_ sensor2_4_ _0372_ _0376_ NAND3
X3787 VSS VDD _0373_ _0374_ _0377_ NOR2
X3788 VSS VDD _0369_ _0372_ _0378_ XOR
X3789 VSS VDD _0368_ _0378_ _0379_ NOR2
X3790 VSS VDD _0355_ _0361_ _0367_ _0379_ _0380_ AOI31
X3791 VSS VDD finestra_gaussiana2_7_ sensor2_5_ _0381_ NAND2
X3792 VSS VDD finestra_gaussiana2_6_ _0366_ _0382_ NAND2
X3793 VSS VDD sensor2_6_ finestra_gaussiana2_6_ _0383_ NAND2
X3794 VSS VDD sensor2_6_ finestra_gaussiana2_6_ _0366_ _0384_ AOI21
X3795 VSS VDD finestra_gaussiana2_6_ _0366_ _0384_ _0385_ AOI21
X3796 VSS VDD _0381_ _0385_ _0387_ XOR
X3797 VSS VDD _0387_ _0388_ INVERTER
X3798 VSS VDD _0365_ _0387_ _0389_ NOR2
X3799 VSS VDD _0365_ _0387_ _0390_ XOR
X3800 VSS VDD _0365_ _0388_ _0391_ XOR
X3801 VSS VDD _0380_ _0391_ _0392_ NOR2
X3802 VSS VDD _0380_ _0390_ _0393_ XOR
X3803 VSS VDD _0369_ _0371_ _0370_ _0394_ OAI21
X3804 VSS VDD _0370_ _0376_ _0393_ _0395_ AOI21
X3805 VSS VDD _0392_ _0395_ _0396_ NOR2
X3806 VSS VDD finestra_gaussiana2_6_ sensor2_7_ _0398_ NAND2
X3807 VSS VDD finestra_gaussiana2_7_ sensor2_6_ _0399_ NAND2
X3808 VSS VDD finestra_gaussiana2_7_ sensor2_7_ _0400_ NAND2
X3809 VSS VDD _0398_ _0399_ _0401_ XOR
X3810 VSS VDD _0389_ _0401_ _0402_ NAND2
X3811 VSS VDD _0389_ _0401_ _0403_ XOR
X3812 VSS VDD _0381_ _0384_ _0382_ _0404_ OAI21
X3813 VSS VDD _0403_ _0404_ _0405_ NAND2
X3814 VSS VDD _0403_ _0404_ _0406_ XOR
X3815 VSS VDD _0392_ _0395_ _0406_ _0407_ OAI21
X3816 VSS VDD _0396_ _0406_ _0409_ XOR
X3817 VSS VDD sensor2_5_ finestra_gaussiana2_3_ _0410_ NAND2
X3818 VSS VDD sensor2_7_ finestra_gaussiana2_1_ _0411_ NAND2
X3819 VSS VDD sensor2_5_ finestra_gaussiana2_1_ _0412_ NAND2
X3820 VSS VDD _0354_ _0412_ _0413_ NOR2
X3821 VSS VDD sensor2_6_ _0413_ _0414_ NAND2
X3822 VSS VDD sensor2_6_ finestra_gaussiana2_3_ _0415_ NAND2
X3823 VSS VDD _0354_ _0412_ _0415_ _0416_ OAI21
X3824 VSS VDD _0414_ _0416_ _0417_ NAND2
X3825 VSS VDD finestra_gaussiana2_5_ sensor2_4_ _0418_ NAND2
X3826 VSS VDD sensor2_7_ finestra_gaussiana2_2_ _0420_ NAND2
X3827 VSS VDD sensor2_5_ finestra_gaussiana2_2_ _0421_ NAND2
X3828 VSS VDD _0363_ _0421_ _0422_ NOR2
X3829 VSS VDD _0359_ _0420_ _0423_ XOR
X3830 VSS VDD _0418_ _0423_ _0424_ XOR
X3831 VSS VDD _0417_ _0424_ _0414_ _0425_ OAI21
X3832 VSS VDD _0355_ _0361_ _0426_ XOR
X3833 VSS VDD _0354_ _0361_ _0427_ XOR
X3834 VSS VDD _0425_ _0427_ _0428_ XOR
X3835 VSS VDD finestra_gaussiana2_7_ sensor2_3_ _0429_ NAND2
X3836 VSS VDD finestra_gaussiana2_6_ sensor2_4_ _0431_ NAND2
X3837 VSS VDD finestra_gaussiana2_5_ sensor2_4_ _0423_ _0422_ _0432_ AOI31
X3838 VSS VDD _0431_ _0432_ _0433_ XOR
X3839 VSS VDD finestra_gaussiana2_7_ sensor2_3_ _0433_ _0434_ NAND3
X3840 VSS VDD _0429_ _0433_ _0435_ XOR
X3841 VSS VDD _0428_ _0435_ _0436_ NOR2
X3842 VSS VDD _0425_ _0426_ _0436_ _0437_ AOI21
X3843 VSS VDD _0368_ _0377_ _0438_ XOR
X3844 VSS VDD _0437_ _0438_ _0439_ NOR2
X3845 VSS VDD _0437_ _0438_ _0440_ XOR
X3846 VSS VDD _0431_ _0432_ _0434_ _0442_ OAI21
X3847 VSS VDD _0440_ _0442_ _0439_ _0443_ AOI21
X3848 VSS VDD _0393_ _0394_ _0444_ XOR
X3849 VSS VDD _0444_ _0445_ INVERTER
X3850 VSS VDD _0443_ _0444_ _0446_ NOR2
X3851 VSS VDD sensor2_7_ finestra_gaussiana2_0_ _0447_ NAND2
X3852 VSS VDD finestra_gaussiana2_3_ sensor2_4_ _0448_ NAND2
X3853 VSS VDD sensor2_4_ finestra_gaussiana2_0_ _0449_ NAND2
X3854 VSS VDD _0354_ _0449_ _0450_ NOR2
X3855 VSS VDD _0447_ _0448_ _0451_ XOR
X3856 VSS VDD sensor2_6_ finestra_gaussiana2_1_ _0453_ NAND2
X3857 VSS VDD sensor2_6_ finestra_gaussiana2_1_ _0451_ _0454_ NAND3
X3858 VSS VDD sensor2_6_ finestra_gaussiana2_1_ _0451_ _0450_ _0455_ AOI31
X3859 VSS VDD _0354_ _0449_ _0454_ _0456_ OAI21
X3860 VSS VDD _0410_ _0411_ _0457_ XOR
X3861 VSS VDD _0456_ _0457_ _0458_ NAND2
X3862 VSS VDD _0455_ _0457_ _0459_ XOR
X3863 VSS VDD finestra_gaussiana2_5_ sensor2_3_ _0460_ NAND2
X3864 VSS VDD finestra_gaussiana2_4_ sensor2_4_ _0461_ NAND2
X3865 VSS VDD sensor2_6_ finestra_gaussiana2_2_ _0462_ NAND2
X3866 VSS VDD sensor2_4_ finestra_gaussiana2_2_ _0464_ NAND2
X3867 VSS VDD _0356_ _0464_ _0465_ NOR2
X3868 VSS VDD _0461_ _0462_ _0466_ XOR
X3869 VSS VDD finestra_gaussiana2_5_ sensor2_3_ _0466_ _0467_ NAND3
X3870 VSS VDD _0460_ _0466_ _0468_ XOR
X3871 VSS VDD _0459_ _0468_ _0469_ NOR2
X3872 VSS VDD _0456_ _0457_ _0469_ _0470_ AOI21
X3873 VSS VDD _0459_ _0468_ _0458_ _0471_ OAI21
X3874 VSS VDD _0417_ _0424_ _0472_ XOR
X3875 VSS VDD _0471_ _0472_ _0473_ NAND2
X3876 VSS VDD _0470_ _0472_ _0475_ XOR
X3877 VSS VDD finestra_gaussiana2_7_ sensor2_2_ _0476_ NAND2
X3878 VSS VDD finestra_gaussiana2_6_ sensor2_3_ _0477_ NAND2
X3879 VSS VDD finestra_gaussiana2_5_ sensor2_3_ _0466_ _0465_ _0478_ AOI31
X3880 VSS VDD _0356_ _0464_ _0467_ _0479_ OAI21
X3881 VSS VDD finestra_gaussiana2_6_ sensor2_3_ _0479_ _0480_ NAND3
X3882 VSS VDD _0477_ _0478_ _0481_ XOR
X3883 VSS VDD finestra_gaussiana2_7_ sensor2_2_ _0481_ _0482_ NAND3
X3884 VSS VDD _0476_ _0481_ _0483_ XOR
X3885 VSS VDD _0475_ _0483_ _0473_ _0484_ OAI21
X3886 VSS VDD _0428_ _0435_ _0486_ XOR
X3887 VSS VDD _0484_ _0486_ _0487_ XOR
X3888 VSS VDD _0487_ _0488_ INVERTER
X3889 VSS VDD _0480_ _0482_ _0489_ NAND2
X3890 VSS VDD _0480_ _0482_ _0488_ _0490_ AOI21
X3891 VSS VDD _0484_ _0486_ _0490_ _0491_ AOI21
X3892 VSS VDD _0491_ _0492_ INVERTER
X3893 VSS VDD _0440_ _0442_ _0493_ XOR
X3894 VSS VDD _0492_ _0493_ _0494_ NAND2
X3895 VSS VDD _0492_ _0493_ _0495_ XOR
X3896 VSS VDD sensor2_6_ finestra_gaussiana2_0_ _0497_ NAND2
X3897 VSS VDD finestra_gaussiana2_3_ sensor2_3_ _0498_ NAND2
X3898 VSS VDD sensor2_3_ finestra_gaussiana2_0_ _0499_ NAND2
X3899 VSS VDD _0415_ _0499_ _0500_ NOR2
X3900 VSS VDD _0497_ _0498_ _0501_ XOR
X3901 VSS VDD sensor2_5_ finestra_gaussiana2_1_ _0501_ _0500_ _0502_ AOI31
X3902 VSS VDD _0451_ _0453_ _0503_ XOR
X3903 VSS VDD _0502_ _0503_ _0504_ XOR
X3904 VSS VDD finestra_gaussiana2_5_ sensor2_2_ _0505_ NAND2
X3905 VSS VDD finestra_gaussiana2_4_ sensor2_3_ _0506_ NAND2
X3906 VSS VDD finestra_gaussiana2_2_ sensor2_3_ _0508_ NAND2
X3907 VSS VDD _0359_ _0508_ _0509_ NOR2
X3908 VSS VDD _0421_ _0506_ _0510_ NAND2
X3909 VSS VDD _0421_ _0506_ _0511_ XOR
X3910 VSS VDD _0359_ _0508_ _0510_ _0512_ OAI21
X3911 VSS VDD finestra_gaussiana2_5_ sensor2_2_ _0511_ _0513_ NAND3
X3912 VSS VDD _0505_ _0512_ _0514_ XOR
X3913 VSS VDD _0505_ _0511_ _0515_ XOR
X3914 VSS VDD _0504_ _0514_ _0516_ NAND2
X3915 VSS VDD _0502_ _0503_ _0516_ _0517_ OAI21
X3916 VSS VDD _0459_ _0468_ _0519_ XOR
X3917 VSS VDD _0517_ _0519_ _0520_ NAND2
X3918 VSS VDD _0517_ _0519_ _0521_ XOR
X3919 VSS VDD finestra_gaussiana2_7_ sensor2_1_ _0522_ NAND2
X3920 VSS VDD finestra_gaussiana2_6_ sensor2_2_ _0523_ NAND2
X3921 VSS VDD finestra_gaussiana2_5_ sensor2_2_ _0510_ _0509_ _0524_ AOI31
X3922 VSS VDD _0359_ _0508_ _0513_ _0525_ OAI21
X3923 VSS VDD finestra_gaussiana2_6_ sensor2_2_ _0525_ _0526_ NAND3
X3924 VSS VDD _0523_ _0524_ _0527_ XOR
X3925 VSS VDD _0523_ _0525_ _0528_ XOR
X3926 VSS VDD finestra_gaussiana2_7_ sensor2_1_ _0527_ _0530_ NAND3
X3927 VSS VDD _0522_ _0528_ _0531_ XOR
X3928 VSS VDD _0521_ _0531_ _0532_ NAND2
X3929 VSS VDD _0520_ _0532_ _0533_ NAND2
X3930 VSS VDD _0533_ _0534_ INVERTER
X3931 VSS VDD _0475_ _0483_ _0535_ XOR
X3932 VSS VDD _0534_ _0535_ _0536_ XOR
X3933 VSS VDD _0526_ _0530_ _0537_ NAND2
X3934 VSS VDD _0526_ _0530_ _0536_ _0538_ AOI21
X3935 VSS VDD _0533_ _0535_ _0538_ _0539_ AOI21
X3936 VSS VDD _0488_ _0489_ _0541_ XOR
X3937 VSS VDD _0541_ _0542_ INVERTER
X3938 VSS VDD _0539_ _0541_ _0543_ NOR2
X3939 VSS VDD _0539_ _0541_ _0544_ XOR
X3940 VSS VDD _0539_ _0542_ _0545_ XOR
X3941 VSS VDD sensor2_5_ finestra_gaussiana2_0_ _0546_ NAND2
X3942 VSS VDD finestra_gaussiana2_3_ sensor2_2_ _0547_ NAND2
X3943 VSS VDD finestra_gaussiana2_0_ sensor2_2_ _0548_ NAND2
X3944 VSS VDD _0546_ _0547_ _0549_ XOR
X3945 VSS VDD sensor2_4_ finestra_gaussiana2_1_ _0550_ NAND2
X3946 VSS VDD sensor2_4_ finestra_gaussiana2_1_ _0549_ _0552_ NAND3
X3947 VSS VDD _0410_ _0548_ _0552_ _0553_ OAI21
X3948 VSS VDD _0412_ _0501_ _0554_ XOR
X3949 VSS VDD _0554_ _0555_ INVERTER
X3950 VSS VDD _0553_ _0555_ _0556_ NAND2
X3951 VSS VDD _0553_ _0554_ _0557_ XOR
X3952 VSS VDD finestra_gaussiana2_5_ sensor2_1_ _0558_ NAND2
X3953 VSS VDD finestra_gaussiana2_4_ sensor2_2_ _0559_ NAND2
X3954 VSS VDD finestra_gaussiana2_2_ sensor2_2_ _0560_ NAND2
X3955 VSS VDD _0464_ _0559_ _0561_ NOR2
X3956 VSS VDD _0464_ _0559_ _0563_ XOR
X3957 VSS VDD _0558_ _0563_ _0564_ XOR
X3958 VSS VDD _0557_ _0564_ _0556_ _0565_ OAI21
X3959 VSS VDD _0504_ _0514_ _0566_ XOR
X3960 VSS VDD _0504_ _0515_ _0567_ XOR
X3961 VSS VDD _0565_ _0566_ _0568_ NAND2
X3962 VSS VDD _0565_ _0567_ _0569_ XOR
X3963 VSS VDD finestra_gaussiana2_7_ sensor2_0_ _0570_ NAND2
X3964 VSS VDD finestra_gaussiana2_6_ sensor2_1_ _0571_ NAND2
X3965 VSS VDD finestra_gaussiana2_5_ sensor2_1_ _0563_ _0561_ _0572_ AOI31
X3966 VSS VDD _0571_ _0572_ _0574_ NOR2
X3967 VSS VDD _0571_ _0572_ _0575_ XOR
X3968 VSS VDD _0570_ _0575_ _0576_ XOR
X3969 VSS VDD _0569_ _0576_ _0568_ _0577_ OAI21
X3970 VSS VDD _0521_ _0531_ _0578_ XOR
X3971 VSS VDD _0577_ _0578_ _0579_ NAND2
X3972 VSS VDD _0577_ _0578_ _0580_ XOR
X3973 VSS VDD _0580_ _0581_ INVERTER
X3974 VSS VDD finestra_gaussiana2_7_ sensor2_0_ _0575_ _0574_ _0582_ AOI31
X3975 VSS VDD _0581_ _0582_ _0583_ NOR2
X3976 VSS VDD _0577_ _0578_ _0583_ _0585_ AOI21
X3977 VSS VDD _0581_ _0582_ _0579_ _0586_ OAI21
X3978 VSS VDD _0536_ _0537_ _0587_ XOR
X3979 VSS VDD _0585_ _0587_ _0588_ NOR2
X3980 VSS VDD _0586_ _0587_ _0589_ XOR
X3981 VSS VDD finestra_gaussiana2_3_ sensor2_1_ _0590_ NAND2
X3982 VSS VDD finestra_gaussiana2_0_ sensor2_1_ _0591_ NAND2
X3983 VSS VDD _0448_ _0591_ _0592_ NOR2
X3984 VSS VDD _0449_ _0590_ _0593_ XOR
X3985 VSS VDD finestra_gaussiana2_1_ sensor2_3_ _0594_ NAND2
X3986 VSS VDD finestra_gaussiana2_1_ sensor2_3_ _0593_ _0592_ _0596_ AOI31
X3987 VSS VDD _0549_ _0550_ _0597_ XOR
X3988 VSS VDD _0596_ _0597_ _0598_ XOR
X3989 VSS VDD finestra_gaussiana2_5_ sensor2_0_ _0599_ NAND2
X3990 VSS VDD finestra_gaussiana2_4_ sensor2_1_ _0600_ NAND2
X3991 VSS VDD finestra_gaussiana2_2_ sensor2_1_ _0601_ NAND2
X3992 VSS VDD _0506_ _0601_ _0602_ NOR2
X3993 VSS VDD _0508_ _0600_ _0603_ NAND2
X3994 VSS VDD _0506_ _0601_ _0603_ _0604_ OAI21
X3995 VSS VDD _0599_ _0604_ _0605_ XOR
X3996 VSS VDD _0598_ _0605_ _0607_ NAND2
X3997 VSS VDD _0596_ _0597_ _0607_ _0608_ OAI21
X3998 VSS VDD _0557_ _0564_ _0609_ XOR
X3999 VSS VDD _0608_ _0609_ _0610_ NAND2
X4000 VSS VDD _0608_ _0609_ _0611_ XOR
X4001 VSS VDD finestra_gaussiana2_6_ sensor2_0_ _0612_ NAND2
X4002 VSS VDD finestra_gaussiana2_5_ sensor2_0_ _0603_ _0602_ _0613_ AOI31
X4003 VSS VDD _0612_ _0613_ _0614_ NOR2
X4004 VSS VDD _0612_ _0613_ _0615_ XOR
X4005 VSS VDD _0611_ _0615_ _0616_ NAND2
X4006 VSS VDD _0610_ _0616_ _0618_ NAND2
X4007 VSS VDD _0569_ _0576_ _0619_ XOR
X4008 VSS VDD _0618_ _0619_ _0620_ NAND2
X4009 VSS VDD _0618_ _0619_ _0621_ XOR
X4010 VSS VDD _0614_ _0621_ _0622_ NAND2
X4011 VSS VDD _0620_ _0622_ _0623_ NAND2
X4012 VSS VDD _0580_ _0582_ _0624_ XOR
X4013 VSS VDD _0620_ _0622_ _0624_ _0625_ AOI21
X4014 VSS VDD _0593_ _0594_ _0626_ XOR
X4015 VSS VDD finestra_gaussiana2_3_ sensor2_0_ _0627_ NAND2
X4016 VSS VDD finestra_gaussiana2_0_ sensor2_0_ _0629_ NAND2
X4017 VSS VDD _0498_ _0629_ _0630_ NOR2
X4018 VSS VDD finestra_gaussiana2_1_ sensor2_2_ _0631_ NAND2
X4019 VSS VDD _0499_ _0627_ _0631_ _0632_ AOI21
X4020 VSS VDD _0630_ _0632_ _0633_ NOR2
X4021 VSS VDD _0626_ _0633_ _0634_ NOR2
X4022 VSS VDD _0626_ _0633_ _0635_ XOR
X4023 VSS VDD finestra_gaussiana2_4_ sensor2_0_ _0636_ NAND2
X4024 VSS VDD finestra_gaussiana2_2_ sensor2_0_ _0637_ NAND2
X4025 VSS VDD _0559_ _0637_ _0638_ NOR2
X4026 VSS VDD _0560_ _0636_ _0640_ XOR
X4027 VSS VDD _0635_ _0640_ _0641_ NAND2
X4028 VSS VDD _0635_ _0640_ _0634_ _0642_ AOI21
X4029 VSS VDD _0626_ _0633_ _0641_ _0643_ OAI21
X4030 VSS VDD _0598_ _0605_ _0644_ XOR
X4031 VSS VDD _0643_ _0644_ _0645_ NAND2
X4032 VSS VDD _0642_ _0644_ _0646_ XOR
X4033 VSS VDD _0646_ _0647_ INVERTER
X4034 VSS VDD _0638_ _0647_ _0648_ NAND2
X4035 VSS VDD _0559_ _0637_ _0645_ _0646_ _0649_ OAI31
X4036 VSS VDD _0611_ _0615_ _0651_ XOR
X4037 VSS VDD _0651_ _0652_ INVERTER
X4038 VSS VDD _0645_ _0648_ _0652_ _0653_ AOI21
X4039 VSS VDD _0649_ _0651_ _0654_ NAND2
X4040 VSS VDD _0614_ _0621_ _0655_ XOR
X4041 VSS VDD _0653_ _0655_ _0656_ NAND2
X4042 VSS VDD _0653_ _0655_ _0657_ XOR
X4043 VSS VDD _0654_ _0655_ _0658_ XOR
X4044 VSS VDD _0499_ _0627_ _0659_ XOR
X4045 VSS VDD finestra_gaussiana2_1_ sensor2_1_ _0660_ NAND2
X4046 VSS VDD _0591_ _0631_ _0659_ _0662_ NOR3
X4047 VSS VDD finestra_gaussiana2_1_ sensor2_2_ _0591_ _0663_ NAND3
X4048 VSS VDD _0659_ _0663_ _0664_ XOR
X4049 VSS VDD _0601_ _0664_ _0665_ NOR2
X4050 VSS VDD _0662_ _0665_ _0666_ NOR2
X4051 VSS VDD _0635_ _0640_ _0667_ XOR
X4052 VSS VDD _0662_ _0665_ _0667_ _0668_ OAI21
X4053 VSS VDD _0638_ _0647_ _0669_ XOR
X4054 VSS VDD _0638_ _0646_ _0670_ XOR
X4055 VSS VDD _0668_ _0670_ _0671_ NOR2
X4056 VSS VDD _0649_ _0651_ _0673_ XOR
X4057 VSS VDD _0671_ _0673_ _0674_ NAND2
X4058 VSS VDD finestra_gaussiana2_1_ sensor2_0_ _0675_ NAND2
X4059 VSS VDD _0629_ _0660_ _0676_ NOR2
X4060 VSS VDD _0548_ _0660_ _0677_ XOR
X4061 VSS VDD _0676_ _0677_ _0678_ NAND2
X4062 VSS VDD _0676_ _0677_ _0679_ NOR2
X4063 VSS VDD _0676_ _0677_ _0680_ XOR
X4064 VSS VDD _0637_ _0679_ _0678_ _0681_ OAI21
X4065 VSS VDD _0601_ _0664_ _0682_ XOR
X4066 VSS VDD _0681_ _0682_ _0684_ NAND2
X4067 VSS VDD _0666_ _0667_ _0685_ XOR
X4068 VSS VDD _0684_ _0685_ _0686_ NOR2
X4069 VSS VDD _0669_ _0686_ _0687_ NAND2
X4070 VSS VDD _0671_ _0673_ _0688_ NOR2
X4071 VSS VDD _0671_ _0673_ _0689_ XOR
X4072 VSS VDD _0687_ _0688_ _0674_ _0690_ OAI21
X4073 VSS VDD _0657_ _0690_ _0691_ NAND2
X4074 VSS VDD _0656_ _0691_ _0692_ NAND2
X4075 VSS VDD _0623_ _0624_ _0693_ XOR
X4076 VSS VDD _0693_ _0695_ INVERTER
X4077 VSS VDD _0692_ _0695_ _0625_ _0696_ AOI21
X4078 VSS VDD _0589_ _0696_ _0697_ NOR2
X4079 VSS VDD _0588_ _0697_ _0698_ NOR2
X4080 VSS VDD _0545_ _0698_ _0699_ NOR2
X4081 VSS VDD _0543_ _0699_ _0700_ NOR2
X4082 VSS VDD _0543_ _0699_ _0495_ _0701_ OAI21
X4083 VSS VDD _0494_ _0701_ _0702_ NAND2
X4084 VSS VDD _0443_ _0445_ _0703_ XOR
X4085 VSS VDD _0703_ _0704_ INVERTER
X4086 VSS VDD _0702_ _0704_ _0446_ _0706_ AOI21
X4087 VSS VDD _0409_ _0706_ _0407_ _0707_ OAI21
X4088 VSS VDD _0402_ _0405_ _0708_ NAND2
X4089 VSS VDD sensor2_6_ finestra_gaussiana2_6_ _0400_ _0709_ AOI21
X4090 VSS VDD finestra_gaussiana2_7_ sensor2_7_ _0383_ _0710_ NAND3
X4091 VSS VDD _0708_ _0709_ _0711_ XOR
X4092 VSS VDD _0708_ _0710_ _0712_ XOR
X4093 VSS VDD _0383_ _0402_ _0405_ _0400_ _0713_ AOI31
X4094 VSS VDD _0707_ _0711_ _0713_ _0714_ AOI21
X4095 VSS VDD sensor3_7_ finestra_gaussiana3_3_ _0715_ NAND2
X4096 VSS VDD _0715_ _0717_ INVERTER
X4097 VSS VDD finestra_gaussiana3_5_ sensor3_5_ _0718_ NAND2
X4098 VSS VDD sensor3_6_ finestra_gaussiana3_4_ _0719_ NAND2
X4099 VSS VDD sensor3_6_ finestra_gaussiana3_5_ _0720_ NAND2
X4100 VSS VDD finestra_gaussiana3_4_ sensor3_5_ _0721_ NAND2
X4101 VSS VDD _0720_ _0721_ _0722_ NOR2
X4102 VSS VDD _0718_ _0719_ _0723_ XOR
X4103 VSS VDD _0717_ _0723_ _0724_ NAND2
X4104 VSS VDD sensor3_7_ finestra_gaussiana3_4_ _0725_ NAND2
X4105 VSS VDD sensor3_7_ finestra_gaussiana3_5_ _0726_ NAND2
X4106 VSS VDD _0719_ _0726_ _0728_ NOR2
X4107 VSS VDD _0720_ _0725_ _0729_ NAND2
X4108 VSS VDD _0720_ _0725_ _0730_ XOR
X4109 VSS VDD _0719_ _0726_ _0729_ _0731_ OAI21
X4110 VSS VDD _0724_ _0731_ _0732_ NOR2
X4111 VSS VDD _0724_ _0731_ _0733_ XOR
X4112 VSS VDD _0724_ _0730_ _0734_ XOR
X4113 VSS VDD finestra_gaussiana3_7_ sensor3_4_ _0735_ NAND2
X4114 VSS VDD finestra_gaussiana3_6_ _0722_ _0736_ NAND2
X4115 VSS VDD finestra_gaussiana3_6_ sensor3_5_ _0722_ _0737_ AOI21
X4116 VSS VDD finestra_gaussiana3_6_ _0722_ _0737_ _0739_ AOI21
X4117 VSS VDD finestra_gaussiana3_6_ _0722_ _0735_ _0737_ _0740_ AOI211
X4118 VSS VDD _0735_ _0739_ _0741_ XOR
X4119 VSS VDD _0734_ _0741_ _0742_ NOR2
X4120 VSS VDD _0732_ _0742_ _0743_ NOR2
X4121 VSS VDD finestra_gaussiana3_7_ sensor3_5_ _0744_ NAND2
X4122 VSS VDD finestra_gaussiana3_6_ _0728_ _0745_ NAND2
X4123 VSS VDD sensor3_6_ finestra_gaussiana3_6_ _0746_ NAND2
X4124 VSS VDD sensor3_6_ finestra_gaussiana3_6_ _0728_ _0747_ AOI21
X4125 VSS VDD finestra_gaussiana3_6_ _0728_ _0747_ _0748_ AOI21
X4126 VSS VDD _0744_ _0748_ _0750_ XOR
X4127 VSS VDD _0726_ _0750_ _0751_ NOR2
X4128 VSS VDD _0726_ _0750_ _0752_ XOR
X4129 VSS VDD _0732_ _0742_ _0752_ _0753_ OAI21
X4130 VSS VDD _0743_ _0752_ _0754_ XOR
X4131 VSS VDD finestra_gaussiana3_6_ _0722_ _0740_ _0755_ AOI21
X4132 VSS VDD _0735_ _0737_ _0736_ _0756_ OAI21
X4133 VSS VDD _0754_ _0755_ _0753_ _0757_ OAI21
X4134 VSS VDD finestra_gaussiana3_6_ sensor3_7_ _0758_ NAND2
X4135 VSS VDD finestra_gaussiana3_7_ sensor3_6_ _0759_ NAND2
X4136 VSS VDD finestra_gaussiana3_7_ sensor3_7_ _0761_ NAND2
X4137 VSS VDD _0758_ _0759_ _0762_ XOR
X4138 VSS VDD _0751_ _0762_ _0763_ NAND2
X4139 VSS VDD _0751_ _0762_ _0764_ XOR
X4140 VSS VDD _0744_ _0747_ _0745_ _0765_ OAI21
X4141 VSS VDD _0764_ _0765_ _0766_ NAND2
X4142 VSS VDD _0764_ _0765_ _0767_ XOR
X4143 VSS VDD _0757_ _0767_ _0768_ NAND2
X4144 VSS VDD _0757_ _0767_ _0769_ XOR
X4145 VSS VDD _0769_ _0770_ INVERTER
X4146 VSS VDD sensor3_5_ finestra_gaussiana3_3_ _0772_ NAND2
X4147 VSS VDD sensor3_7_ finestra_gaussiana3_1_ _0773_ NAND2
X4148 VSS VDD sensor3_5_ finestra_gaussiana3_1_ _0774_ NAND2
X4149 VSS VDD _0715_ _0774_ _0775_ NOR2
X4150 VSS VDD sensor3_6_ _0775_ _0776_ NAND2
X4151 VSS VDD sensor3_6_ finestra_gaussiana3_3_ _0777_ NAND2
X4152 VSS VDD _0715_ _0774_ _0777_ _0778_ OAI21
X4153 VSS VDD _0776_ _0778_ _0779_ NAND2
X4154 VSS VDD finestra_gaussiana3_5_ sensor3_4_ _0780_ NAND2
X4155 VSS VDD sensor3_7_ finestra_gaussiana3_2_ _0781_ NAND2
X4156 VSS VDD sensor3_5_ finestra_gaussiana3_2_ _0783_ NAND2
X4157 VSS VDD _0725_ _0783_ _0784_ NOR2
X4158 VSS VDD _0721_ _0781_ _0785_ XOR
X4159 VSS VDD _0780_ _0785_ _0786_ XOR
X4160 VSS VDD _0779_ _0786_ _0776_ _0787_ OAI21
X4161 VSS VDD _0717_ _0723_ _0788_ XOR
X4162 VSS VDD _0715_ _0723_ _0789_ XOR
X4163 VSS VDD _0787_ _0789_ _0790_ XOR
X4164 VSS VDD finestra_gaussiana3_7_ sensor3_3_ _0791_ NAND2
X4165 VSS VDD finestra_gaussiana3_6_ sensor3_4_ _0792_ NAND2
X4166 VSS VDD finestra_gaussiana3_5_ sensor3_4_ _0785_ _0784_ _0794_ AOI31
X4167 VSS VDD _0792_ _0794_ _0795_ XOR
X4168 VSS VDD finestra_gaussiana3_7_ sensor3_3_ _0795_ _0796_ NAND3
X4169 VSS VDD _0791_ _0795_ _0797_ XOR
X4170 VSS VDD _0790_ _0797_ _0798_ NOR2
X4171 VSS VDD _0787_ _0788_ _0798_ _0799_ AOI21
X4172 VSS VDD _0733_ _0741_ _0800_ XOR
X4173 VSS VDD _0799_ _0800_ _0801_ NOR2
X4174 VSS VDD _0799_ _0800_ _0802_ XOR
X4175 VSS VDD _0792_ _0794_ _0796_ _0803_ OAI21
X4176 VSS VDD _0802_ _0803_ _0801_ _0805_ AOI21
X4177 VSS VDD _0754_ _0756_ _0806_ XOR
X4178 VSS VDD _0806_ _0807_ INVERTER
X4179 VSS VDD _0805_ _0806_ _0808_ NOR2
X4180 VSS VDD sensor3_7_ finestra_gaussiana3_0_ _0809_ NAND2
X4181 VSS VDD finestra_gaussiana3_3_ sensor3_4_ _0810_ NAND2
X4182 VSS VDD sensor3_4_ finestra_gaussiana3_0_ _0811_ NAND2
X4183 VSS VDD _0715_ _0811_ _0812_ NOR2
X4184 VSS VDD _0809_ _0810_ _0813_ XOR
X4185 VSS VDD sensor3_6_ finestra_gaussiana3_1_ _0814_ NAND2
X4186 VSS VDD sensor3_6_ finestra_gaussiana3_1_ _0813_ _0816_ NAND3
X4187 VSS VDD sensor3_6_ finestra_gaussiana3_1_ _0813_ _0812_ _0817_ AOI31
X4188 VSS VDD _0715_ _0811_ _0816_ _0818_ OAI21
X4189 VSS VDD _0772_ _0773_ _0819_ XOR
X4190 VSS VDD _0818_ _0819_ _0820_ NAND2
X4191 VSS VDD _0817_ _0819_ _0821_ XOR
X4192 VSS VDD finestra_gaussiana3_5_ sensor3_3_ _0822_ NAND2
X4193 VSS VDD finestra_gaussiana3_4_ sensor3_4_ _0823_ NAND2
X4194 VSS VDD sensor3_6_ finestra_gaussiana3_2_ _0824_ NAND2
X4195 VSS VDD sensor3_4_ finestra_gaussiana3_2_ _0825_ NAND2
X4196 VSS VDD _0719_ _0825_ _0827_ NOR2
X4197 VSS VDD _0823_ _0824_ _0828_ XOR
X4198 VSS VDD finestra_gaussiana3_5_ sensor3_3_ _0828_ _0829_ NAND3
X4199 VSS VDD _0822_ _0828_ _0830_ XOR
X4200 VSS VDD _0821_ _0830_ _0831_ NOR2
X4201 VSS VDD _0818_ _0819_ _0831_ _0832_ AOI21
X4202 VSS VDD _0821_ _0830_ _0820_ _0833_ OAI21
X4203 VSS VDD _0779_ _0786_ _0834_ XOR
X4204 VSS VDD _0833_ _0834_ _0835_ NAND2
X4205 VSS VDD _0832_ _0834_ _0836_ XOR
X4206 VSS VDD finestra_gaussiana3_7_ sensor3_2_ _0838_ NAND2
X4207 VSS VDD finestra_gaussiana3_6_ sensor3_3_ _0839_ NAND2
X4208 VSS VDD finestra_gaussiana3_5_ sensor3_3_ _0828_ _0827_ _0840_ AOI31
X4209 VSS VDD _0719_ _0825_ _0829_ _0841_ OAI21
X4210 VSS VDD finestra_gaussiana3_6_ sensor3_3_ _0841_ _0842_ NAND3
X4211 VSS VDD _0839_ _0840_ _0843_ XOR
X4212 VSS VDD finestra_gaussiana3_7_ sensor3_2_ _0843_ _0844_ NAND3
X4213 VSS VDD _0838_ _0843_ _0845_ XOR
X4214 VSS VDD _0836_ _0845_ _0835_ _0846_ OAI21
X4215 VSS VDD _0790_ _0797_ _0847_ XOR
X4216 VSS VDD _0846_ _0847_ _0849_ XOR
X4217 VSS VDD _0849_ _0850_ INVERTER
X4218 VSS VDD _0842_ _0844_ _0851_ NAND2
X4219 VSS VDD _0842_ _0844_ _0850_ _0852_ AOI21
X4220 VSS VDD _0846_ _0847_ _0852_ _0853_ AOI21
X4221 VSS VDD _0853_ _0854_ INVERTER
X4222 VSS VDD _0802_ _0803_ _0855_ XOR
X4223 VSS VDD _0854_ _0855_ _0856_ NAND2
X4224 VSS VDD _0853_ _0855_ _0857_ XOR
X4225 VSS VDD _0857_ _0858_ INVERTER
X4226 VSS VDD sensor3_6_ finestra_gaussiana3_0_ _0860_ NAND2
X4227 VSS VDD finestra_gaussiana3_3_ sensor3_3_ _0861_ NAND2
X4228 VSS VDD sensor3_3_ finestra_gaussiana3_0_ _0862_ NAND2
X4229 VSS VDD _0777_ _0862_ _0863_ NOR2
X4230 VSS VDD _0860_ _0861_ _0864_ XOR
X4231 VSS VDD sensor3_5_ finestra_gaussiana3_1_ _0864_ _0863_ _0865_ AOI31
X4232 VSS VDD _0813_ _0814_ _0866_ XOR
X4233 VSS VDD _0865_ _0866_ _0867_ XOR
X4234 VSS VDD finestra_gaussiana3_5_ sensor3_2_ _0868_ NAND2
X4235 VSS VDD finestra_gaussiana3_4_ sensor3_3_ _0869_ NAND2
X4236 VSS VDD finestra_gaussiana3_2_ sensor3_3_ _0871_ NAND2
X4237 VSS VDD _0783_ _0869_ _0872_ NAND2
X4238 VSS VDD _0783_ _0869_ _0873_ XOR
X4239 VSS VDD _0721_ _0871_ _0872_ _0874_ OAI21
X4240 VSS VDD finestra_gaussiana3_5_ sensor3_2_ _0873_ _0875_ NAND3
X4241 VSS VDD _0868_ _0874_ _0876_ XOR
X4242 VSS VDD _0868_ _0873_ _0877_ XOR
X4243 VSS VDD _0867_ _0876_ _0878_ NAND2
X4244 VSS VDD _0865_ _0866_ _0878_ _0879_ OAI21
X4245 VSS VDD _0821_ _0830_ _0880_ XOR
X4246 VSS VDD _0879_ _0880_ _0882_ NAND2
X4247 VSS VDD _0879_ _0880_ _0883_ XOR
X4248 VSS VDD finestra_gaussiana3_7_ sensor3_1_ _0884_ NAND2
X4249 VSS VDD finestra_gaussiana3_6_ sensor3_2_ _0885_ NAND2
X4250 VSS VDD _0721_ _0871_ _0875_ _0886_ OAI21
X4251 VSS VDD finestra_gaussiana3_6_ sensor3_2_ _0886_ _0887_ NAND3
X4252 VSS VDD _0885_ _0886_ _0888_ XOR
X4253 VSS VDD _0884_ _0888_ _0889_ XOR
X4254 VSS VDD _0883_ _0889_ _0890_ NAND2
X4255 VSS VDD _0882_ _0890_ _0891_ NAND2
X4256 VSS VDD _0836_ _0845_ _0893_ XOR
X4257 VSS VDD _0891_ _0893_ _0894_ NAND2
X4258 VSS VDD _0891_ _0893_ _0895_ XOR
X4259 VSS VDD _0884_ _0888_ _0887_ _0896_ OAI21
X4260 VSS VDD _0896_ _0897_ INVERTER
X4261 VSS VDD _0895_ _0896_ _0898_ NAND2
X4262 VSS VDD _0894_ _0898_ _0899_ NAND2
X4263 VSS VDD _0850_ _0851_ _0900_ XOR
X4264 VSS VDD _0894_ _0898_ _0900_ _0901_ AOI21
X4265 VSS VDD _0899_ _0900_ _0902_ XOR
X4266 VSS VDD _0902_ _0904_ INVERTER
X4267 VSS VDD sensor3_5_ finestra_gaussiana3_0_ _0905_ NAND2
X4268 VSS VDD finestra_gaussiana3_3_ sensor3_2_ _0906_ NAND2
X4269 VSS VDD finestra_gaussiana3_0_ sensor3_2_ _0907_ NAND2
X4270 VSS VDD _0905_ _0906_ _0908_ XOR
X4271 VSS VDD sensor3_4_ finestra_gaussiana3_1_ _0909_ NAND2
X4272 VSS VDD sensor3_4_ finestra_gaussiana3_1_ _0908_ _0910_ NAND3
X4273 VSS VDD _0772_ _0907_ _0910_ _0911_ OAI21
X4274 VSS VDD _0774_ _0864_ _0912_ XOR
X4275 VSS VDD _0912_ _0913_ INVERTER
X4276 VSS VDD _0911_ _0913_ _0915_ NAND2
X4277 VSS VDD _0911_ _0912_ _0916_ XOR
X4278 VSS VDD finestra_gaussiana3_5_ sensor3_1_ _0917_ NAND2
X4279 VSS VDD finestra_gaussiana3_4_ sensor3_2_ _0918_ NAND2
X4280 VSS VDD finestra_gaussiana3_2_ sensor3_2_ _0919_ NAND2
X4281 VSS VDD _0825_ _0918_ _0920_ NOR2
X4282 VSS VDD _0825_ _0918_ _0921_ XOR
X4283 VSS VDD _0917_ _0921_ _0922_ XOR
X4284 VSS VDD _0916_ _0922_ _0915_ _0923_ OAI21
X4285 VSS VDD _0867_ _0876_ _0924_ XOR
X4286 VSS VDD _0867_ _0877_ _0926_ XOR
X4287 VSS VDD _0923_ _0924_ _0927_ NAND2
X4288 VSS VDD _0923_ _0926_ _0928_ XOR
X4289 VSS VDD finestra_gaussiana3_7_ sensor3_0_ _0929_ NAND2
X4290 VSS VDD finestra_gaussiana3_6_ sensor3_1_ _0930_ NAND2
X4291 VSS VDD finestra_gaussiana3_5_ sensor3_1_ _0921_ _0920_ _0931_ AOI31
X4292 VSS VDD _0930_ _0931_ _0932_ NOR2
X4293 VSS VDD _0930_ _0931_ _0933_ XOR
X4294 VSS VDD _0929_ _0933_ _0934_ XOR
X4295 VSS VDD _0928_ _0934_ _0927_ _0935_ OAI21
X4296 VSS VDD _0883_ _0889_ _0937_ XOR
X4297 VSS VDD _0935_ _0937_ _0938_ XOR
X4298 VSS VDD _0938_ _0939_ INVERTER
X4299 VSS VDD finestra_gaussiana3_7_ sensor3_0_ _0933_ _0932_ _0940_ AOI31
X4300 VSS VDD _0939_ _0940_ _0941_ NOR2
X4301 VSS VDD _0935_ _0937_ _0941_ _0942_ AOI21
X4302 VSS VDD _0895_ _0896_ _0943_ XOR
X4303 VSS VDD _0895_ _0897_ _0944_ XOR
X4304 VSS VDD _0942_ _0944_ _0945_ NOR2
X4305 VSS VDD _0942_ _0943_ _0946_ XOR
X4306 VSS VDD _0946_ _0948_ INVERTER
X4307 VSS VDD finestra_gaussiana3_3_ sensor3_1_ _0949_ NAND2
X4308 VSS VDD finestra_gaussiana3_0_ sensor3_1_ _0950_ NAND2
X4309 VSS VDD _0810_ _0950_ _0951_ NOR2
X4310 VSS VDD _0811_ _0949_ _0952_ XOR
X4311 VSS VDD finestra_gaussiana3_1_ sensor3_3_ _0953_ NAND2
X4312 VSS VDD finestra_gaussiana3_1_ sensor3_3_ _0952_ _0951_ _0954_ AOI31
X4313 VSS VDD _0908_ _0909_ _0955_ XOR
X4314 VSS VDD _0954_ _0955_ _0956_ XOR
X4315 VSS VDD finestra_gaussiana3_5_ sensor3_0_ _0957_ NAND2
X4316 VSS VDD finestra_gaussiana3_4_ sensor3_1_ _0959_ NAND2
X4317 VSS VDD finestra_gaussiana3_2_ sensor3_1_ _0960_ NAND2
X4318 VSS VDD _0869_ _0960_ _0961_ NOR2
X4319 VSS VDD _0871_ _0959_ _0962_ NAND2
X4320 VSS VDD _0869_ _0960_ _0962_ _0963_ OAI21
X4321 VSS VDD _0957_ _0963_ _0964_ XOR
X4322 VSS VDD _0956_ _0964_ _0965_ NAND2
X4323 VSS VDD _0954_ _0955_ _0965_ _0966_ OAI21
X4324 VSS VDD _0916_ _0922_ _0967_ XOR
X4325 VSS VDD _0966_ _0967_ _0968_ NAND2
X4326 VSS VDD _0966_ _0967_ _0970_ XOR
X4327 VSS VDD finestra_gaussiana3_6_ sensor3_0_ _0971_ NAND2
X4328 VSS VDD finestra_gaussiana3_5_ sensor3_0_ _0962_ _0961_ _0972_ AOI31
X4329 VSS VDD _0971_ _0972_ _0973_ NOR2
X4330 VSS VDD _0971_ _0972_ _0974_ XOR
X4331 VSS VDD _0970_ _0974_ _0975_ NAND2
X4332 VSS VDD _0968_ _0975_ _0976_ NAND2
X4333 VSS VDD _0928_ _0934_ _0977_ XOR
X4334 VSS VDD _0976_ _0977_ _0978_ NAND2
X4335 VSS VDD _0976_ _0977_ _0979_ NOR2
X4336 VSS VDD _0976_ _0977_ _0981_ XOR
X4337 VSS VDD _0971_ _0972_ _0978_ _0979_ _0982_ OAI31
X4338 VSS VDD _0939_ _0940_ _0983_ XOR
X4339 VSS VDD _0982_ _0983_ _0984_ NAND2
X4340 VSS VDD _0952_ _0953_ _0985_ XOR
X4341 VSS VDD finestra_gaussiana3_3_ sensor3_0_ _0986_ NAND2
X4342 VSS VDD finestra_gaussiana3_0_ sensor3_0_ _0987_ NAND2
X4343 VSS VDD _0861_ _0987_ _0988_ NOR2
X4344 VSS VDD finestra_gaussiana3_1_ sensor3_2_ _0989_ NAND2
X4345 VSS VDD _0862_ _0986_ _0989_ _0990_ AOI21
X4346 VSS VDD _0988_ _0990_ _0992_ NOR2
X4347 VSS VDD _0985_ _0992_ _0993_ NOR2
X4348 VSS VDD _0985_ _0992_ _0994_ XOR
X4349 VSS VDD finestra_gaussiana3_4_ sensor3_0_ _0995_ NAND2
X4350 VSS VDD finestra_gaussiana3_2_ sensor3_0_ _0996_ NAND2
X4351 VSS VDD _0918_ _0996_ _0997_ NOR2
X4352 VSS VDD _0919_ _0995_ _0998_ XOR
X4353 VSS VDD _0994_ _0998_ _0999_ NAND2
X4354 VSS VDD _0994_ _0998_ _0993_ _1000_ AOI21
X4355 VSS VDD _0985_ _0992_ _0999_ _1001_ OAI21
X4356 VSS VDD _0956_ _0964_ _1003_ XOR
X4357 VSS VDD _1001_ _1003_ _1004_ NAND2
X4358 VSS VDD _1000_ _1003_ _1005_ XOR
X4359 VSS VDD _0918_ _0996_ _1004_ _1005_ _1006_ OAI31
X4360 VSS VDD _0970_ _0974_ _1007_ XOR
X4361 VSS VDD _1006_ _1007_ _1008_ NAND2
X4362 VSS VDD _0973_ _0981_ _1009_ XOR
X4363 VSS VDD _1009_ _1010_ INVERTER
X4364 VSS VDD _1008_ _1010_ _1011_ NOR2
X4365 VSS VDD _0862_ _0986_ _1012_ XOR
X4366 VSS VDD finestra_gaussiana3_1_ sensor3_1_ _1014_ NAND2
X4367 VSS VDD _0950_ _0989_ _1012_ _1015_ NOR3
X4368 VSS VDD finestra_gaussiana3_0_ sensor3_1_ _0989_ _1016_ AOI21
X4369 VSS VDD finestra_gaussiana3_1_ sensor3_2_ _0950_ _1017_ NAND3
X4370 VSS VDD _1012_ _1017_ _1018_ XOR
X4371 VSS VDD _1012_ _1016_ _1019_ XOR
X4372 VSS VDD finestra_gaussiana3_2_ sensor3_1_ _1019_ _1020_ NAND3
X4373 VSS VDD finestra_gaussiana3_2_ sensor3_1_ _1019_ _1015_ _1021_ AOI31
X4374 VSS VDD _0950_ _0989_ _1020_ _1012_ _1022_ OAI31
X4375 VSS VDD _0994_ _0998_ _1023_ XOR
X4376 VSS VDD _1022_ _1023_ _1025_ NAND2
X4377 VSS VDD _0997_ _1005_ _1026_ XOR
X4378 VSS VDD _1025_ _1026_ _1027_ NOR2
X4379 VSS VDD _1006_ _1007_ _1028_ XOR
X4380 VSS VDD _1027_ _1028_ _1029_ NAND2
X4381 VSS VDD finestra_gaussiana3_1_ sensor3_0_ _1030_ NAND2
X4382 VSS VDD _0987_ _1014_ _1031_ NOR2
X4383 VSS VDD _0907_ _1014_ _1032_ XOR
X4384 VSS VDD finestra_gaussiana3_0_ sensor3_2_ _0987_ _1014_ _1033_ AOI211
X4385 VSS VDD _1031_ _1032_ _1034_ NOR2
X4386 VSS VDD _1031_ _1032_ _1036_ XOR
X4387 VSS VDD _0996_ _1033_ _1034_ _1037_ NOR3
X4388 VSS VDD finestra_gaussiana3_2_ sensor3_0_ _1036_ _1033_ _1038_ AOI31
X4389 VSS VDD _0960_ _1018_ _1039_ XOR
X4390 VSS VDD _1033_ _1037_ _1039_ _1040_ OAI21
X4391 VSS VDD _1022_ _1023_ _1041_ XOR
X4392 VSS VDD _1021_ _1023_ _1042_ XOR
X4393 VSS VDD _1026_ _1040_ _1042_ _1043_ NOR3
X4394 VSS VDD _1043_ _1044_ INVERTER
X4395 VSS VDD _1027_ _1028_ _1045_ XOR
X4396 VSS VDD _1043_ _1045_ _1047_ NAND2
X4397 VSS VDD _1029_ _1047_ _1048_ NAND2
X4398 VSS VDD _1008_ _1010_ _1049_ XOR
X4399 VSS VDD _1008_ _1009_ _1050_ XOR
X4400 VSS VDD _1029_ _1047_ _1050_ _1051_ AOI21
X4401 VSS VDD _1011_ _1051_ _1052_ NOR2
X4402 VSS VDD _0982_ _0983_ _1053_ XOR
X4403 VSS VDD _1011_ _1051_ _1053_ _1054_ OAI21
X4404 VSS VDD _0984_ _1054_ _1055_ NAND2
X4405 VSS VDD _0948_ _1055_ _0945_ _1056_ AOI21
X4406 VSS VDD _0902_ _1056_ _1058_ NOR2
X4407 VSS VDD _0901_ _1058_ _1059_ NOR2
X4408 VSS VDD _0901_ _1058_ _0858_ _1060_ OAI21
X4409 VSS VDD _0856_ _1060_ _1061_ NAND2
X4410 VSS VDD _0805_ _0807_ _1062_ XOR
X4411 VSS VDD _0856_ _1060_ _1062_ _1063_ AOI21
X4412 VSS VDD _0808_ _1063_ _1064_ NOR2
X4413 VSS VDD _0770_ _1064_ _0768_ _1065_ OAI21
X4414 VSS VDD _0763_ _0766_ _1066_ NAND2
X4415 VSS VDD sensor3_6_ finestra_gaussiana3_6_ _0761_ _1067_ AOI21
X4416 VSS VDD _1066_ _1067_ _1069_ NAND2
X4417 VSS VDD _1066_ _1067_ _1070_ XOR
X4418 VSS VDD _1070_ _1071_ INVERTER
X4419 VSS VDD _1065_ _1070_ _1072_ NAND2
X4420 VSS VDD _1065_ _1071_ _1073_ XOR
X4421 VSS VDD _0341_ _0344_ _1074_ XOR
X4422 VSS VDD _1073_ _1074_ _1075_ NOR2
X4423 VSS VDD _0770_ _1064_ _1076_ XOR
X4424 VSS VDD _0769_ _1064_ _1077_ XOR
X4425 VSS VDD _0252_ _0340_ _1078_ XOR
X4426 VSS VDD _1076_ _1078_ _1080_ NAND2
X4427 VSS VDD _1076_ _1078_ _1081_ XOR
X4428 VSS VDD _1077_ _1078_ _1082_ XOR
X4429 VSS VDD _1061_ _1062_ _1083_ XOR
X4430 VSS VDD _0258_ _0339_ _1084_ XOR
X4431 VSS VDD _1083_ _1084_ _1085_ NOR2
X4432 VSS VDD _0857_ _1059_ _1086_ XOR
X4433 VSS VDD _0259_ _0260_ _1087_ XOR
X4434 VSS VDD _0259_ _0261_ _1088_ XOR
X4435 VSS VDD _0338_ _1087_ _1089_ XOR
X4436 VSS VDD _0338_ _1088_ _1091_ XOR
X4437 VSS VDD _1086_ _1091_ _1092_ NAND2
X4438 VSS VDD _1086_ _1091_ _1093_ XOR
X4439 VSS VDD _1086_ _1089_ _1094_ XOR
X4440 VSS VDD _0904_ _1056_ _1095_ XOR
X4441 VSS VDD _0267_ _0337_ _1096_ XOR
X4442 VSS VDD _1095_ _1096_ _1097_ NOR2
X4443 VSS VDD _1095_ _1096_ _1098_ XOR
X4444 VSS VDD _0948_ _1055_ _1099_ XOR
X4445 VSS VDD _0946_ _1055_ _1100_ XOR
X4446 VSS VDD _0268_ _0270_ _1102_ XOR
X4447 VSS VDD _0335_ _1102_ _1103_ XOR
X4448 VSS VDD _1099_ _1103_ _1104_ NAND2
X4449 VSS VDD _1099_ _1103_ _1105_ XOR
X4450 VSS VDD _1100_ _1103_ _1106_ XOR
X4451 VSS VDD _1052_ _1053_ _1107_ XOR
X4452 VSS VDD _0332_ _0333_ _1108_ XOR
X4453 VSS VDD _1107_ _1108_ _1109_ NOR2
X4454 VSS VDD _1048_ _1049_ _1110_ XOR
X4455 VSS VDD _1048_ _1050_ _1111_ XOR
X4456 VSS VDD _0282_ _0330_ _1113_ XOR
X4457 VSS VDD _1110_ _1113_ _1114_ NAND2
X4458 VSS VDD _1110_ _1113_ _1115_ XOR
X4459 VSS VDD _1111_ _1113_ _1116_ XOR
X4460 VSS VDD _1044_ _1045_ _1117_ XOR
X4461 VSS VDD _0288_ _0329_ _1118_ XOR
X4462 VSS VDD _1117_ _1118_ _1119_ NOR2
X4463 VSS VDD _1117_ _1118_ _1120_ XOR
X4464 VSS VDD _0295_ _0328_ _1121_ XOR
X4465 VSS VDD _1040_ _1042_ _1025_ _1122_ OAI21
X4466 VSS VDD _1026_ _1122_ _1124_ XOR
X4467 VSS VDD _1124_ _1125_ INVERTER
X4468 VSS VDD _1121_ _1125_ _1126_ NAND2
X4469 VSS VDD _1121_ _1125_ _1127_ XOR
X4470 VSS VDD _1121_ _1124_ _1128_ XOR
X4471 VSS VDD _1040_ _1042_ _1129_ XOR
X4472 VSS VDD _1040_ _1041_ _1130_ XOR
X4473 VSS VDD _0324_ _0326_ _1131_ XOR
X4474 VSS VDD _1130_ _1131_ _1132_ NOR2
X4475 VSS VDD _1038_ _1039_ _1133_ XOR
X4476 VSS VDD _0303_ _0322_ _1135_ XOR
X4477 VSS VDD _1133_ _1135_ _1136_ NOR2
X4478 VSS VDD _1133_ _1135_ _1137_ XOR
X4479 VSS VDD _0996_ _1036_ _1138_ XOR
X4480 VSS VDD _0317_ _0318_ _1139_ XOR
X4481 VSS VDD _0317_ _0319_ _1140_ XOR
X4482 VSS VDD _1138_ _1140_ _1141_ NOR2
X4483 VSS VDD _0950_ _1030_ _1142_ XOR
X4484 VSS VDD _0314_ _0316_ _1143_ XOR
X4485 VSS VDD _1142_ _1143_ _1144_ NAND2
X4486 VSS VDD _1928_ _0312_ _1146_ XOR
X4487 VSS VDD _0987_ _1146_ _1147_ NOR2
X4488 VSS VDD _1142_ _1143_ _1148_ NOR2
X4489 VSS VDD _1142_ _1143_ _1149_ XOR
X4490 VSS VDD _0987_ _1148_ _1144_ _1146_ _1150_ OAI31
X4491 VSS VDD _1138_ _1140_ _1151_ XOR
X4492 VSS VDD _1138_ _1139_ _1152_ XOR
X4493 VSS VDD _1150_ _1151_ _1153_ NAND2
X4494 VSS VDD _1150_ _1151_ _1141_ _1154_ AOI21
X4495 VSS VDD _1138_ _1140_ _1153_ _1155_ OAI21
X4496 VSS VDD _1137_ _1155_ _1136_ _1157_ AOI21
X4497 VSS VDD _1130_ _1131_ _1158_ XOR
X4498 VSS VDD _1129_ _1131_ _1159_ XOR
X4499 VSS VDD _1157_ _1159_ _1160_ NOR2
X4500 VSS VDD _1132_ _1160_ _1161_ NOR2
X4501 VSS VDD _1128_ _1161_ _1126_ _1162_ OAI21
X4502 VSS VDD _1120_ _1162_ _1119_ _1163_ AOI21
X4503 VSS VDD _1116_ _1163_ _1114_ _1164_ OAI21
X4504 VSS VDD _1107_ _1108_ _1165_ XOR
X4505 VSS VDD _1164_ _1165_ _1109_ _1166_ AOI21
X4506 VSS VDD _1106_ _1166_ _1104_ _1168_ OAI21
X4507 VSS VDD _1098_ _1168_ _1097_ _1169_ AOI21
X4508 VSS VDD _1094_ _1169_ _1092_ _1170_ OAI21
X4509 VSS VDD _1083_ _1084_ _1171_ XOR
X4510 VSS VDD _1170_ _1171_ _1085_ _1172_ AOI21
X4511 VSS VDD _1082_ _1172_ _1080_ _1173_ OAI21
X4512 VSS VDD _1073_ _1074_ _1174_ XOR
X4513 VSS VDD _1173_ _1174_ _1075_ _1175_ AOI21
X4514 VSS VDD _0746_ _0763_ _0766_ _0761_ _1176_ AOI31
X4515 VSS VDD _1065_ _1070_ _1176_ _1177_ AOI21
X4516 VSS VDD _0746_ _0761_ _1069_ _1072_ _1179_ OAI211
X4517 VSS VDD _0345_ _0346_ _1180_ XOR
X4518 VSS VDD _1180_ _1181_ INVERTER
X4519 VSS VDD _1177_ _1180_ _1182_ XOR
X4520 VSS VDD _1179_ _1180_ _1183_ XOR
X4521 VSS VDD _1175_ _1183_ _1184_ NOR2
X4522 VSS VDD _1175_ _1183_ _1185_ XOR
X4523 VSS VDD _1175_ _1182_ _1186_ XOR
X4524 VSS VDD _0714_ _1186_ _1187_ NOR2
X4525 VSS VDD _0714_ _1186_ _1188_ XOR
X4526 VSS VDD _0714_ _1185_ _1190_ XOR
X4527 VSS VDD _0707_ _0711_ _1191_ XOR
X4528 VSS VDD _0707_ _0712_ _1192_ XOR
X4529 VSS VDD _1173_ _1174_ _1193_ XOR
X4530 VSS VDD _1191_ _1193_ _1194_ NAND2
X4531 VSS VDD _1191_ _1193_ _1195_ XOR
X4532 VSS VDD _1192_ _1193_ _1196_ XOR
X4533 VSS VDD _0409_ _0706_ _1197_ XOR
X4534 VSS VDD _1197_ _1198_ INVERTER
X4535 VSS VDD _1082_ _1172_ _1199_ XOR
X4536 VSS VDD _1081_ _1172_ _1201_ XOR
X4537 VSS VDD _1198_ _1201_ _1202_ NOR2
X4538 VSS VDD _1197_ _1199_ _1203_ XOR
X4539 VSS VDD _1198_ _1199_ _1204_ XOR
X4540 VSS VDD _0702_ _0704_ _1205_ XOR
X4541 VSS VDD _0702_ _0703_ _1206_ XOR
X4542 VSS VDD _1170_ _1171_ _1207_ XOR
X4543 VSS VDD _1205_ _1207_ _1208_ NAND2
X4544 VSS VDD _1205_ _1207_ _1209_ XOR
X4545 VSS VDD _1206_ _1207_ _1210_ XOR
X4546 VSS VDD _0495_ _0700_ _1212_ XOR
X4547 VSS VDD _1094_ _1169_ _1213_ XOR
X4548 VSS VDD _1093_ _1169_ _1214_ XOR
X4549 VSS VDD _1212_ _1214_ _1215_ NOR2
X4550 VSS VDD _1212_ _1214_ _1216_ XOR
X4551 VSS VDD _1212_ _1213_ _1217_ XOR
X4552 VSS VDD _0545_ _0698_ _1218_ XOR
X4553 VSS VDD _0544_ _0698_ _1219_ XOR
X4554 VSS VDD _1098_ _1168_ _1220_ XOR
X4555 VSS VDD _1218_ _1220_ _1221_ NAND2
X4556 VSS VDD _1219_ _1220_ _1223_ XOR
X4557 VSS VDD _0589_ _0696_ _1224_ XOR
X4558 VSS VDD _1224_ _1225_ INVERTER
X4559 VSS VDD _1106_ _1166_ _1226_ XOR
X4560 VSS VDD _1105_ _1166_ _1227_ XOR
X4561 VSS VDD _1225_ _1227_ _1228_ NOR2
X4562 VSS VDD _1224_ _1226_ _1229_ XOR
X4563 VSS VDD _1225_ _1226_ _1230_ XOR
X4564 VSS VDD _0692_ _0695_ _1231_ XOR
X4565 VSS VDD _0692_ _0693_ _1232_ XOR
X4566 VSS VDD _1164_ _1165_ _1234_ XOR
X4567 VSS VDD _1231_ _1234_ _1235_ NAND2
X4568 VSS VDD _0658_ _0690_ _1236_ XOR
X4569 VSS VDD _1116_ _1163_ _1237_ XOR
X4570 VSS VDD _1115_ _1163_ _1238_ XOR
X4571 VSS VDD _1236_ _1238_ _1239_ NOR2
X4572 VSS VDD _1236_ _1238_ _1240_ XOR
X4573 VSS VDD _1236_ _1237_ _1241_ XOR
X4574 VSS VDD _0687_ _0689_ _1242_ XOR
X4575 VSS VDD _1242_ _1243_ INVERTER
X4576 VSS VDD _1120_ _1162_ _1245_ XOR
X4577 VSS VDD _1243_ _1245_ _1246_ NAND2
X4578 VSS VDD _1242_ _1245_ _1247_ XOR
X4579 VSS VDD _0684_ _0685_ _0668_ _1248_ OAI21
X4580 VSS VDD _0670_ _1248_ _1249_ XOR
X4581 VSS VDD _1127_ _1161_ _1250_ XOR
X4582 VSS VDD _1249_ _1250_ _1251_ NOR2
X4583 VSS VDD _1249_ _1250_ _1252_ XOR
X4584 VSS VDD _0684_ _0685_ _1253_ XOR
X4585 VSS VDD _1157_ _1158_ _1254_ XOR
X4586 VSS VDD _1254_ _1256_ INVERTER
X4587 VSS VDD _1253_ _1256_ _1257_ NAND2
X4588 VSS VDD _0681_ _0682_ _1258_ XOR
X4589 VSS VDD _1137_ _1155_ _1259_ XOR
X4590 VSS VDD _1137_ _1154_ _1260_ XOR
X4591 VSS VDD _1258_ _1260_ _1261_ XOR
X4592 VSS VDD _0637_ _0680_ _1262_ XOR
X4593 VSS VDD _1150_ _1151_ _1263_ XOR
X4594 VSS VDD _1150_ _1152_ _1264_ XOR
X4595 VSS VDD _1262_ _1264_ _1265_ NOR2
X4596 VSS VDD _0591_ _0675_ _1267_ XOR
X4597 VSS VDD _1147_ _1149_ _1268_ XOR
X4598 VSS VDD _1267_ _1268_ _1269_ NAND2
X4599 VSS VDD _0987_ _1146_ _1270_ XOR
X4600 VSS VDD _1270_ _1271_ INVERTER
X4601 VSS VDD _0629_ _1271_ _1272_ NOR2
X4602 VSS VDD _1267_ _1268_ _1273_ NOR2
X4603 VSS VDD _1267_ _1268_ _1274_ XOR
X4604 VSS VDD _0629_ _1273_ _1269_ _1271_ _1275_ OAI31
X4605 VSS VDD _1262_ _1264_ _1276_ XOR
X4606 VSS VDD _1262_ _1263_ _1278_ XOR
X4607 VSS VDD _1275_ _1276_ _1265_ _1279_ AOI21
X4608 VSS VDD _1261_ _1279_ _1280_ NOR2
X4609 VSS VDD _1258_ _1259_ _1280_ _1281_ AOI21
X4610 VSS VDD _1253_ _1254_ _1282_ XOR
X4611 VSS VDD _1281_ _1282_ _1283_ NOR2
X4612 VSS VDD _1253_ _1256_ _1283_ _1284_ AOI21
X4613 VSS VDD _1281_ _1282_ _1257_ _1285_ OAI21
X4614 VSS VDD _1252_ _1285_ _1251_ _1286_ AOI21
X4615 VSS VDD _1247_ _1286_ _1246_ _1287_ OAI21
X4616 VSS VDD _1240_ _1287_ _1239_ _1289_ AOI21
X4617 VSS VDD _1232_ _1234_ _1290_ XOR
X4618 VSS VDD _1289_ _1290_ _1235_ _1291_ OAI21
X4619 VSS VDD _1229_ _1291_ _1228_ _1292_ AOI21
X4620 VSS VDD _1223_ _1292_ _1221_ _1293_ OAI21
X4621 VSS VDD _1216_ _1293_ _1215_ _1294_ AOI21
X4622 VSS VDD _1210_ _1294_ _1208_ _1295_ OAI21
X4623 VSS VDD _1203_ _1295_ _1202_ _1296_ AOI21
X4624 VSS VDD _1196_ _1296_ _1194_ _1297_ OAI21
X4625 VSS VDD _1188_ _1297_ _1187_ _1298_ AOI21
X4626 VSS VDD _1179_ _1181_ _1184_ _1300_ AOI21
X4627 VSS VDD _0349_ _0350_ _1301_ XOR
X4628 VSS VDD _0349_ _0351_ _1302_ XOR
X4629 VSS VDD _1300_ _1302_ _1303_ NOR2
X4630 VSS VDD _1300_ _1302_ _1304_ XOR
X4631 VSS VDD _1300_ _1301_ _1305_ XOR
X4632 VSS VDD _1298_ _1305_ _1306_ NOR2
X4633 VSS VDD _0349_ _0350_ _1298_ _1300_ _1307_ NOR4
X4634 VSS VDD _0352_ _1306_ _1308_ NAND2
X4635 VSS VDD _0352_ _1303_ _1309_ NOR2
X4636 VSS VDD _0352_ _1303_ _1306_ _1311_ NOR3
X4637 VSS VDD _1298_ _1305_ _1309_ _1312_ OAI21
X4638 VSS VDD sensor1_7_ finestra_gaussiana1_3_ _1313_ NAND2
X4639 VSS VDD _1313_ _1314_ INVERTER
X4640 VSS VDD sensor1_6_ finestra_gaussiana1_4_ _1315_ NAND2
X4641 VSS VDD finestra_gaussiana1_5_ sensor1_5_ _1316_ NAND2
X4642 VSS VDD sensor1_6_ finestra_gaussiana1_5_ _1317_ NAND2
X4643 VSS VDD finestra_gaussiana1_4_ sensor1_5_ _1318_ NAND2
X4644 VSS VDD _1317_ _1318_ _1319_ NOR2
X4645 VSS VDD _1315_ _1316_ _1320_ XOR
X4646 VSS VDD _1314_ _1320_ _1322_ NAND2
X4647 VSS VDD sensor1_7_ finestra_gaussiana1_4_ _1323_ NAND2
X4648 VSS VDD sensor1_7_ finestra_gaussiana1_5_ _1324_ NAND2
X4649 VSS VDD _1315_ _1324_ _1325_ NOR2
X4650 VSS VDD _1317_ _1323_ _1326_ NAND2
X4651 VSS VDD _1317_ _1323_ _1327_ XOR
X4652 VSS VDD _1315_ _1324_ _1326_ _1328_ OAI21
X4653 VSS VDD _1322_ _1328_ _1329_ NOR2
X4654 VSS VDD _1322_ _1328_ _1330_ XOR
X4655 VSS VDD _1322_ _1327_ _1331_ XOR
X4656 VSS VDD finestra_gaussiana1_7_ sensor1_4_ _1333_ NAND2
X4657 VSS VDD finestra_gaussiana1_6_ _1319_ _1334_ NAND2
X4658 VSS VDD finestra_gaussiana1_6_ sensor1_5_ _1319_ _1335_ AOI21
X4659 VSS VDD finestra_gaussiana1_6_ _1319_ _1335_ _1336_ AOI21
X4660 VSS VDD finestra_gaussiana1_6_ _1319_ _1333_ _1335_ _1337_ AOI211
X4661 VSS VDD _1333_ _1336_ _1338_ XOR
X4662 VSS VDD _1331_ _1338_ _1339_ NOR2
X4663 VSS VDD _1329_ _1339_ _1340_ NOR2
X4664 VSS VDD finestra_gaussiana1_7_ sensor1_5_ _1341_ NAND2
X4665 VSS VDD finestra_gaussiana1_6_ _1325_ _1342_ NAND2
X4666 VSS VDD sensor1_6_ finestra_gaussiana1_6_ _1344_ NAND2
X4667 VSS VDD sensor1_6_ finestra_gaussiana1_6_ _1325_ _1345_ AOI21
X4668 VSS VDD finestra_gaussiana1_6_ _1325_ _1345_ _1346_ AOI21
X4669 VSS VDD _1341_ _1346_ _1347_ XOR
X4670 VSS VDD _1324_ _1347_ _1348_ NOR2
X4671 VSS VDD _1324_ _1347_ _1349_ XOR
X4672 VSS VDD _1329_ _1339_ _1349_ _1350_ OAI21
X4673 VSS VDD _1340_ _1349_ _1351_ XOR
X4674 VSS VDD finestra_gaussiana1_6_ _1319_ _1337_ _1352_ AOI21
X4675 VSS VDD _1333_ _1335_ _1334_ _1353_ OAI21
X4676 VSS VDD _1351_ _1352_ _1350_ _1355_ OAI21
X4677 VSS VDD finestra_gaussiana1_6_ sensor1_7_ _1356_ NAND2
X4678 VSS VDD finestra_gaussiana1_7_ sensor1_6_ _1357_ NAND2
X4679 VSS VDD finestra_gaussiana1_7_ sensor1_7_ _1358_ NAND2
X4680 VSS VDD _1356_ _1357_ _1359_ XOR
X4681 VSS VDD _1348_ _1359_ _1360_ NAND2
X4682 VSS VDD _1348_ _1359_ _1361_ XOR
X4683 VSS VDD _1341_ _1345_ _1342_ _1362_ OAI21
X4684 VSS VDD _1361_ _1362_ _1363_ NAND2
X4685 VSS VDD _1361_ _1362_ _1364_ XOR
X4686 VSS VDD _1355_ _1364_ _1366_ NAND2
X4687 VSS VDD _1355_ _1364_ _1367_ XOR
X4688 VSS VDD _1367_ _1368_ INVERTER
X4689 VSS VDD sensor1_5_ finestra_gaussiana1_3_ _1369_ NAND2
X4690 VSS VDD sensor1_7_ finestra_gaussiana1_1_ _1370_ NAND2
X4691 VSS VDD sensor1_5_ finestra_gaussiana1_1_ _1371_ NAND2
X4692 VSS VDD _1313_ _1371_ _1372_ NOR2
X4693 VSS VDD sensor1_6_ _1372_ _1373_ NAND2
X4694 VSS VDD sensor1_6_ finestra_gaussiana1_3_ _1374_ NAND2
X4695 VSS VDD _1313_ _1371_ _1374_ _1375_ OAI21
X4696 VSS VDD _1373_ _1375_ _1377_ NAND2
X4697 VSS VDD finestra_gaussiana1_5_ sensor1_4_ _1378_ NAND2
X4698 VSS VDD sensor1_7_ finestra_gaussiana1_2_ _1379_ NAND2
X4699 VSS VDD sensor1_5_ finestra_gaussiana1_2_ _1380_ NAND2
X4700 VSS VDD _1323_ _1380_ _1381_ NOR2
X4701 VSS VDD _1318_ _1379_ _1382_ XOR
X4702 VSS VDD _1378_ _1382_ _1383_ XOR
X4703 VSS VDD _1377_ _1383_ _1373_ _1384_ OAI21
X4704 VSS VDD _1314_ _1320_ _1385_ XOR
X4705 VSS VDD _1313_ _1320_ _1386_ XOR
X4706 VSS VDD _1384_ _1386_ _1388_ XOR
X4707 VSS VDD finestra_gaussiana1_7_ sensor1_3_ _1389_ NAND2
X4708 VSS VDD finestra_gaussiana1_6_ sensor1_4_ _1390_ NAND2
X4709 VSS VDD finestra_gaussiana1_5_ sensor1_4_ _1382_ _1381_ _1391_ AOI31
X4710 VSS VDD _1390_ _1391_ _1392_ XOR
X4711 VSS VDD finestra_gaussiana1_7_ sensor1_3_ _1392_ _1393_ NAND3
X4712 VSS VDD _1389_ _1392_ _1394_ XOR
X4713 VSS VDD _1388_ _1394_ _1395_ NOR2
X4714 VSS VDD _1384_ _1385_ _1395_ _1396_ AOI21
X4715 VSS VDD _1330_ _1338_ _1397_ XOR
X4716 VSS VDD _1396_ _1397_ _1399_ NOR2
X4717 VSS VDD _1396_ _1397_ _1400_ XOR
X4718 VSS VDD _1390_ _1391_ _1393_ _1401_ OAI21
X4719 VSS VDD _1400_ _1401_ _1399_ _1402_ AOI21
X4720 VSS VDD _1351_ _1353_ _1403_ XOR
X4721 VSS VDD _1402_ _1403_ _1404_ NOR2
X4722 VSS VDD sensor1_7_ finestra_gaussiana1_0_ _1405_ NAND2
X4723 VSS VDD finestra_gaussiana1_3_ sensor1_4_ _1406_ NAND2
X4724 VSS VDD sensor1_4_ finestra_gaussiana1_0_ _1407_ NAND2
X4725 VSS VDD _1313_ _1407_ _1408_ NOR2
X4726 VSS VDD _1405_ _1406_ _1410_ XOR
X4727 VSS VDD sensor1_6_ finestra_gaussiana1_1_ _1411_ NAND2
X4728 VSS VDD sensor1_6_ finestra_gaussiana1_1_ _1410_ _1412_ NAND3
X4729 VSS VDD sensor1_6_ finestra_gaussiana1_1_ _1410_ _1408_ _1413_ AOI31
X4730 VSS VDD _1313_ _1407_ _1412_ _1414_ OAI21
X4731 VSS VDD _1369_ _1370_ _1415_ XOR
X4732 VSS VDD _1414_ _1415_ _1416_ NAND2
X4733 VSS VDD _1413_ _1415_ _1417_ XOR
X4734 VSS VDD finestra_gaussiana1_5_ sensor1_3_ _1418_ NAND2
X4735 VSS VDD finestra_gaussiana1_4_ sensor1_4_ _1419_ NAND2
X4736 VSS VDD sensor1_6_ finestra_gaussiana1_2_ _1421_ NAND2
X4737 VSS VDD sensor1_4_ finestra_gaussiana1_2_ _1422_ NAND2
X4738 VSS VDD _1315_ _1422_ _1423_ NOR2
X4739 VSS VDD _1419_ _1421_ _1424_ XOR
X4740 VSS VDD finestra_gaussiana1_5_ sensor1_3_ _1424_ _1425_ NAND3
X4741 VSS VDD _1418_ _1424_ _1426_ XOR
X4742 VSS VDD _1417_ _1426_ _1427_ NOR2
X4743 VSS VDD _1414_ _1415_ _1427_ _1428_ AOI21
X4744 VSS VDD _1417_ _1426_ _1416_ _1429_ OAI21
X4745 VSS VDD _1377_ _1383_ _1430_ XOR
X4746 VSS VDD _1429_ _1430_ _1432_ NAND2
X4747 VSS VDD _1428_ _1430_ _1433_ XOR
X4748 VSS VDD finestra_gaussiana1_7_ sensor1_2_ _1434_ NAND2
X4749 VSS VDD finestra_gaussiana1_6_ sensor1_3_ _1435_ NAND2
X4750 VSS VDD finestra_gaussiana1_5_ sensor1_3_ _1424_ _1423_ _1436_ AOI31
X4751 VSS VDD _1315_ _1422_ _1425_ _1437_ OAI21
X4752 VSS VDD finestra_gaussiana1_6_ sensor1_3_ _1437_ _1438_ NAND3
X4753 VSS VDD _1435_ _1436_ _1439_ XOR
X4754 VSS VDD finestra_gaussiana1_7_ sensor1_2_ _1439_ _1440_ NAND3
X4755 VSS VDD _1434_ _1439_ _1441_ XOR
X4756 VSS VDD _1433_ _1441_ _1432_ _1443_ OAI21
X4757 VSS VDD _1388_ _1394_ _1444_ XOR
X4758 VSS VDD _1443_ _1444_ _1445_ XOR
X4759 VSS VDD _1445_ _1446_ INVERTER
X4760 VSS VDD _1438_ _1440_ _1447_ NAND2
X4761 VSS VDD _1438_ _1440_ _1446_ _1448_ AOI21
X4762 VSS VDD _1443_ _1444_ _1448_ _1449_ AOI21
X4763 VSS VDD _1449_ _1450_ INVERTER
X4764 VSS VDD _1400_ _1401_ _1451_ XOR
X4765 VSS VDD _1450_ _1451_ _1452_ NAND2
X4766 VSS VDD _1450_ _1451_ _1454_ XOR
X4767 VSS VDD _1449_ _1451_ _1455_ XOR
X4768 VSS VDD sensor1_6_ finestra_gaussiana1_0_ _1456_ NAND2
X4769 VSS VDD finestra_gaussiana1_3_ sensor1_3_ _1457_ NAND2
X4770 VSS VDD sensor1_3_ finestra_gaussiana1_0_ _1458_ NAND2
X4771 VSS VDD _1374_ _1458_ _1459_ NOR2
X4772 VSS VDD _1456_ _1457_ _1460_ XOR
X4773 VSS VDD sensor1_5_ finestra_gaussiana1_1_ _1460_ _1459_ _1461_ AOI31
X4774 VSS VDD _1410_ _1411_ _1462_ XOR
X4775 VSS VDD _1461_ _1462_ _1463_ XOR
X4776 VSS VDD finestra_gaussiana1_5_ sensor1_2_ _1465_ NAND2
X4777 VSS VDD finestra_gaussiana1_4_ sensor1_3_ _1466_ NAND2
X4778 VSS VDD finestra_gaussiana1_2_ sensor1_3_ _1467_ NAND2
X4779 VSS VDD _1318_ _1467_ _1468_ NOR2
X4780 VSS VDD _1380_ _1466_ _1469_ NAND2
X4781 VSS VDD _1380_ _1466_ _1470_ XOR
X4782 VSS VDD _1318_ _1467_ _1469_ _1471_ OAI21
X4783 VSS VDD finestra_gaussiana1_5_ sensor1_2_ _1470_ _1472_ NAND3
X4784 VSS VDD _1465_ _1471_ _1473_ XOR
X4785 VSS VDD _1465_ _1470_ _1474_ XOR
X4786 VSS VDD _1463_ _1473_ _1476_ NAND2
X4787 VSS VDD _1461_ _1462_ _1476_ _1477_ OAI21
X4788 VSS VDD _1417_ _1426_ _1478_ XOR
X4789 VSS VDD _1477_ _1478_ _1479_ NAND2
X4790 VSS VDD _1477_ _1478_ _1480_ XOR
X4791 VSS VDD finestra_gaussiana1_7_ sensor1_1_ _1481_ NAND2
X4792 VSS VDD finestra_gaussiana1_6_ sensor1_2_ _1482_ NAND2
X4793 VSS VDD finestra_gaussiana1_5_ sensor1_2_ _1469_ _1468_ _1483_ AOI31
X4794 VSS VDD _1318_ _1467_ _1472_ _1484_ OAI21
X4795 VSS VDD finestra_gaussiana1_6_ sensor1_2_ _1484_ _1485_ NAND3
X4796 VSS VDD _1482_ _1483_ _1487_ XOR
X4797 VSS VDD _1482_ _1484_ _1488_ XOR
X4798 VSS VDD finestra_gaussiana1_7_ sensor1_1_ _1487_ _1489_ NAND3
X4799 VSS VDD _1481_ _1488_ _1490_ XOR
X4800 VSS VDD _1480_ _1490_ _1491_ NAND2
X4801 VSS VDD _1479_ _1491_ _1492_ NAND2
X4802 VSS VDD _1492_ _1493_ INVERTER
X4803 VSS VDD _1433_ _1441_ _1494_ XOR
X4804 VSS VDD _1493_ _1494_ _1495_ XOR
X4805 VSS VDD _1485_ _1489_ _1496_ NAND2
X4806 VSS VDD _1485_ _1489_ _1495_ _1498_ AOI21
X4807 VSS VDD _1492_ _1494_ _1498_ _1499_ AOI21
X4808 VSS VDD _1446_ _1447_ _1500_ XOR
X4809 VSS VDD _1500_ _1501_ INVERTER
X4810 VSS VDD _1499_ _1500_ _1502_ NOR2
X4811 VSS VDD _1499_ _1501_ _1503_ XOR
X4812 VSS VDD sensor1_5_ finestra_gaussiana1_0_ _1504_ NAND2
X4813 VSS VDD finestra_gaussiana1_3_ sensor1_2_ _1505_ NAND2
X4814 VSS VDD finestra_gaussiana1_0_ sensor1_2_ _1506_ NAND2
X4815 VSS VDD _1504_ _1505_ _1507_ XOR
X4816 VSS VDD sensor1_4_ finestra_gaussiana1_1_ _1509_ NAND2
X4817 VSS VDD sensor1_4_ finestra_gaussiana1_1_ _1507_ _1510_ NAND3
X4818 VSS VDD _1369_ _1506_ _1510_ _1511_ OAI21
X4819 VSS VDD _1371_ _1460_ _1512_ XOR
X4820 VSS VDD _1512_ _1513_ INVERTER
X4821 VSS VDD _1511_ _1513_ _1514_ NAND2
X4822 VSS VDD _1511_ _1512_ _1515_ XOR
X4823 VSS VDD finestra_gaussiana1_5_ sensor1_1_ _1516_ NAND2
X4824 VSS VDD finestra_gaussiana1_4_ sensor1_2_ _1517_ NAND2
X4825 VSS VDD finestra_gaussiana1_2_ sensor1_2_ _1518_ NAND2
X4826 VSS VDD _1422_ _1517_ _1520_ NOR2
X4827 VSS VDD _1422_ _1517_ _1521_ XOR
X4828 VSS VDD _1516_ _1521_ _1522_ XOR
X4829 VSS VDD _1515_ _1522_ _1514_ _1523_ OAI21
X4830 VSS VDD _1463_ _1473_ _1524_ XOR
X4831 VSS VDD _1463_ _1474_ _1525_ XOR
X4832 VSS VDD _1523_ _1524_ _1526_ NAND2
X4833 VSS VDD _1523_ _1525_ _1527_ XOR
X4834 VSS VDD finestra_gaussiana1_7_ sensor1_0_ _1528_ NAND2
X4835 VSS VDD finestra_gaussiana1_6_ sensor1_1_ _1529_ NAND2
X4836 VSS VDD finestra_gaussiana1_5_ sensor1_1_ _1521_ _1520_ _1531_ AOI31
X4837 VSS VDD _1529_ _1531_ _1532_ NOR2
X4838 VSS VDD _1529_ _1531_ _1533_ XOR
X4839 VSS VDD _1528_ _1533_ _1534_ XOR
X4840 VSS VDD _1527_ _1534_ _1526_ _1535_ OAI21
X4841 VSS VDD _1480_ _1490_ _1536_ XOR
X4842 VSS VDD _1535_ _1536_ _1537_ NAND2
X4843 VSS VDD _1535_ _1536_ _1538_ XOR
X4844 VSS VDD _1538_ _1539_ INVERTER
X4845 VSS VDD finestra_gaussiana1_7_ sensor1_0_ _1533_ _1532_ _1540_ AOI31
X4846 VSS VDD _1539_ _1540_ _1542_ NOR2
X4847 VSS VDD _1535_ _1536_ _1542_ _1543_ AOI21
X4848 VSS VDD _1539_ _1540_ _1537_ _1544_ OAI21
X4849 VSS VDD _1495_ _1496_ _1545_ XOR
X4850 VSS VDD _1543_ _1545_ _1546_ NOR2
X4851 VSS VDD _1544_ _1545_ _1547_ XOR
X4852 VSS VDD _1547_ _1548_ INVERTER
X4853 VSS VDD finestra_gaussiana1_3_ sensor1_1_ _1549_ NAND2
X4854 VSS VDD finestra_gaussiana1_0_ sensor1_1_ _1550_ NAND2
X4855 VSS VDD _1406_ _1550_ _1551_ NOR2
X4856 VSS VDD _1407_ _1549_ _1553_ XOR
X4857 VSS VDD finestra_gaussiana1_1_ sensor1_3_ _1554_ NAND2
X4858 VSS VDD finestra_gaussiana1_1_ sensor1_3_ _1553_ _1551_ _1555_ AOI31
X4859 VSS VDD _1507_ _1509_ _1556_ XOR
X4860 VSS VDD _1555_ _1556_ _1557_ XOR
X4861 VSS VDD finestra_gaussiana1_5_ sensor1_0_ _1558_ NAND2
X4862 VSS VDD finestra_gaussiana1_4_ sensor1_1_ _1559_ NAND2
X4863 VSS VDD finestra_gaussiana1_2_ sensor1_1_ _1560_ NAND2
X4864 VSS VDD _1466_ _1560_ _1561_ NOR2
X4865 VSS VDD _1467_ _1559_ _1562_ NAND2
X4866 VSS VDD _1466_ _1560_ _1562_ _1564_ OAI21
X4867 VSS VDD _1558_ _1564_ _1565_ XOR
X4868 VSS VDD _1557_ _1565_ _1566_ NAND2
X4869 VSS VDD _1555_ _1556_ _1566_ _1567_ OAI21
X4870 VSS VDD _1515_ _1522_ _1568_ XOR
X4871 VSS VDD _1567_ _1568_ _1569_ NAND2
X4872 VSS VDD _1567_ _1568_ _1570_ XOR
X4873 VSS VDD finestra_gaussiana1_6_ sensor1_0_ _1571_ NAND2
X4874 VSS VDD finestra_gaussiana1_5_ sensor1_0_ _1562_ _1561_ _1572_ AOI31
X4875 VSS VDD _1571_ _1572_ _1573_ NOR2
X4876 VSS VDD _1571_ _1572_ _1575_ XOR
X4877 VSS VDD _1570_ _1575_ _1576_ NAND2
X4878 VSS VDD _1569_ _1576_ _1577_ NAND2
X4879 VSS VDD _1527_ _1534_ _1578_ XOR
X4880 VSS VDD _1577_ _1578_ _1579_ NAND2
X4881 VSS VDD _1577_ _1578_ _1580_ XOR
X4882 VSS VDD _1573_ _1580_ _1581_ NAND2
X4883 VSS VDD _1579_ _1581_ _1582_ NAND2
X4884 VSS VDD _1538_ _1540_ _1583_ XOR
X4885 VSS VDD _1579_ _1581_ _1583_ _1584_ AOI21
X4886 VSS VDD _1553_ _1554_ _1586_ XOR
X4887 VSS VDD finestra_gaussiana1_3_ sensor1_0_ _1587_ NAND2
X4888 VSS VDD _1458_ _1587_ _1588_ NAND2
X4889 VSS VDD finestra_gaussiana1_0_ sensor1_0_ _1589_ NAND2
X4890 VSS VDD _1457_ _1589_ _1590_ NOR2
X4891 VSS VDD finestra_gaussiana1_1_ sensor1_2_ _1588_ _1590_ _1591_ AOI31
X4892 VSS VDD _1586_ _1591_ _1592_ NOR2
X4893 VSS VDD _1586_ _1591_ _1593_ XOR
X4894 VSS VDD finestra_gaussiana1_4_ sensor1_0_ _1594_ NAND2
X4895 VSS VDD finestra_gaussiana1_2_ sensor1_0_ _1595_ NAND2
X4896 VSS VDD _1517_ _1595_ _1597_ NOR2
X4897 VSS VDD _1518_ _1594_ _1598_ XOR
X4898 VSS VDD _1593_ _1598_ _1599_ NAND2
X4899 VSS VDD _1593_ _1598_ _1592_ _1600_ AOI21
X4900 VSS VDD _1586_ _1591_ _1599_ _1601_ OAI21
X4901 VSS VDD _1557_ _1565_ _1602_ XOR
X4902 VSS VDD _1601_ _1602_ _1603_ NAND2
X4903 VSS VDD _1600_ _1602_ _1604_ XOR
X4904 VSS VDD _1604_ _1605_ INVERTER
X4905 VSS VDD _1597_ _1605_ _1606_ NAND2
X4906 VSS VDD _1517_ _1595_ _1603_ _1604_ _1608_ OAI31
X4907 VSS VDD _1570_ _1575_ _1609_ XOR
X4908 VSS VDD _1609_ _1610_ INVERTER
X4909 VSS VDD _1603_ _1606_ _1610_ _1611_ AOI21
X4910 VSS VDD _1608_ _1609_ _1612_ NAND2
X4911 VSS VDD _1573_ _1580_ _1613_ XOR
X4912 VSS VDD _1611_ _1613_ _1614_ NAND2
X4913 VSS VDD _1611_ _1613_ _1615_ XOR
X4914 VSS VDD _1612_ _1613_ _1616_ XOR
X4915 VSS VDD _1458_ _1587_ _1617_ XOR
X4916 VSS VDD finestra_gaussiana1_1_ sensor1_1_ _1619_ NAND2
X4917 VSS VDD _1506_ _1617_ _1619_ _1620_ NOR3
X4918 VSS VDD finestra_gaussiana1_1_ sensor1_2_ _1550_ _1621_ NAND3
X4919 VSS VDD _1617_ _1621_ _1622_ XOR
X4920 VSS VDD _1560_ _1622_ _1623_ NOR2
X4921 VSS VDD _1620_ _1623_ _1624_ NOR2
X4922 VSS VDD _1593_ _1598_ _1625_ XOR
X4923 VSS VDD _1620_ _1623_ _1625_ _1626_ OAI21
X4924 VSS VDD _1597_ _1605_ _1627_ XOR
X4925 VSS VDD _1597_ _1604_ _1628_ XOR
X4926 VSS VDD _1626_ _1628_ _1630_ NOR2
X4927 VSS VDD _1608_ _1609_ _1631_ XOR
X4928 VSS VDD _1630_ _1631_ _1632_ NAND2
X4929 VSS VDD finestra_gaussiana1_1_ sensor1_0_ _1633_ NAND2
X4930 VSS VDD _1589_ _1619_ _1634_ NOR2
X4931 VSS VDD _1506_ _1619_ _1635_ XOR
X4932 VSS VDD _1634_ _1635_ _1636_ NAND2
X4933 VSS VDD _1634_ _1635_ _1637_ NOR2
X4934 VSS VDD _1634_ _1635_ _1638_ XOR
X4935 VSS VDD _1595_ _1637_ _1636_ _1639_ OAI21
X4936 VSS VDD _1560_ _1622_ _1641_ XOR
X4937 VSS VDD _1639_ _1641_ _1642_ NAND2
X4938 VSS VDD _1624_ _1625_ _1643_ XOR
X4939 VSS VDD _1643_ _1644_ INVERTER
X4940 VSS VDD _1642_ _1643_ _1645_ NOR2
X4941 VSS VDD _1627_ _1645_ _1646_ NAND2
X4942 VSS VDD _1630_ _1631_ _1647_ NOR2
X4943 VSS VDD _1630_ _1631_ _1648_ XOR
X4944 VSS VDD _1646_ _1647_ _1632_ _1649_ OAI21
X4945 VSS VDD _1615_ _1649_ _1650_ NAND2
X4946 VSS VDD _1614_ _1650_ _1652_ NAND2
X4947 VSS VDD _1582_ _1583_ _1653_ XOR
X4948 VSS VDD _1653_ _1654_ INVERTER
X4949 VSS VDD _1652_ _1654_ _1584_ _1655_ AOI21
X4950 VSS VDD _1547_ _1655_ _1656_ NOR2
X4951 VSS VDD _1546_ _1656_ _1657_ NOR2
X4952 VSS VDD _1503_ _1657_ _1658_ NOR2
X4953 VSS VDD _1502_ _1658_ _1659_ NOR2
X4954 VSS VDD _1455_ _1659_ _1452_ _1660_ OAI21
X4955 VSS VDD _1660_ _1661_ INVERTER
X4956 VSS VDD _1402_ _1403_ _1663_ XOR
X4957 VSS VDD _1660_ _1663_ _1404_ _1664_ AOI21
X4958 VSS VDD _1368_ _1664_ _1366_ _1665_ OAI21
X4959 VSS VDD _1360_ _1363_ _1666_ NAND2
X4960 VSS VDD sensor1_6_ finestra_gaussiana1_6_ _1358_ _1667_ AOI21
X4961 VSS VDD finestra_gaussiana1_7_ sensor1_7_ _1344_ _1668_ NAND3
X4962 VSS VDD _1666_ _1667_ _1669_ NAND2
X4963 VSS VDD _1666_ _1667_ _1670_ XOR
X4964 VSS VDD _1666_ _1668_ _1671_ XOR
X4965 VSS VDD _1665_ _1670_ _1672_ NAND2
X4966 VSS VDD _1344_ _1358_ _1669_ _1672_ _1674_ OAI211
X4967 VSS VDD _1674_ _1675_ INVERTER
X4968 VSS VDD _1188_ _1297_ _1676_ XOR
X4969 VSS VDD _1190_ _1297_ _1677_ XOR
X4970 VSS VDD _1675_ _1677_ _1678_ NOR2
X4971 VSS VDD _1674_ _1676_ _1679_ NAND2
X4972 VSS VDD _1674_ _1676_ _1680_ XOR
X4973 VSS VDD _1675_ _1676_ _1681_ XOR
X4974 VSS VDD _1665_ _1670_ _1682_ XOR
X4975 VSS VDD _1665_ _1671_ _1683_ XOR
X4976 VSS VDD _1196_ _1296_ _1685_ XOR
X4977 VSS VDD _1195_ _1296_ _1686_ XOR
X4978 VSS VDD _1683_ _1686_ _1687_ NOR2
X4979 VSS VDD _1682_ _1685_ _1688_ NAND2
X4980 VSS VDD _1682_ _1685_ _1689_ XOR
X4981 VSS VDD _1683_ _1685_ _1690_ XOR
X4982 VSS VDD _1368_ _1664_ _1691_ XOR
X4983 VSS VDD _1367_ _1664_ _1692_ XOR
X4984 VSS VDD _1203_ _1295_ _1693_ XOR
X4985 VSS VDD _1204_ _1295_ _1694_ XOR
X4986 VSS VDD _1692_ _1694_ _1696_ NOR2
X4987 VSS VDD _1691_ _1693_ _1697_ NAND2
X4988 VSS VDD _1691_ _1693_ _1698_ XOR
X4989 VSS VDD _1692_ _1693_ _1699_ XOR
X4990 VSS VDD _1660_ _1663_ _1700_ XOR
X4991 VSS VDD _1661_ _1663_ _1701_ XOR
X4992 VSS VDD _1210_ _1294_ _1702_ XOR
X4993 VSS VDD _1209_ _1294_ _1703_ XOR
X4994 VSS VDD _1700_ _1702_ _1704_ NOR2
X4995 VSS VDD _1701_ _1703_ _1705_ NOR2
X4996 VSS VDD _1700_ _1702_ _1707_ NAND2
X4997 VSS VDD _1455_ _1659_ _1708_ XOR
X4998 VSS VDD _1454_ _1659_ _1709_ XOR
X4999 VSS VDD _1216_ _1293_ _1710_ XOR
X5000 VSS VDD _1217_ _1293_ _1711_ XOR
X5001 VSS VDD _1708_ _1710_ _1712_ NOR2
X5002 VSS VDD _1709_ _1711_ _1713_ NAND2
X5003 VSS VDD _1709_ _1711_ _1714_ NOR2
X5004 VSS VDD _1503_ _1657_ _1715_ XOR
X5005 VSS VDD _1223_ _1292_ _1716_ XOR
X5006 VSS VDD _1715_ _1716_ _1718_ NOR2
X5007 VSS VDD _1715_ _1716_ _1719_ NAND2
X5008 VSS VDD _1548_ _1655_ _1720_ XOR
X5009 VSS VDD _1230_ _1291_ _1721_ XOR
X5010 VSS VDD _1720_ _1721_ _1722_ NOR2
X5011 VSS VDD _1720_ _1721_ _1723_ NAND2
X5012 VSS VDD _1652_ _1654_ _1724_ XOR
X5013 VSS VDD _1289_ _1290_ _1725_ XOR
X5014 VSS VDD _1724_ _1725_ _1726_ NAND2
X5015 VSS VDD _1724_ _1725_ _1727_ NOR2
X5016 VSS VDD _1616_ _1649_ _1729_ XOR
X5017 VSS VDD _1241_ _1287_ _1730_ XOR
X5018 VSS VDD _1729_ _1730_ _1731_ NOR2
X5019 VSS VDD _1729_ _1730_ _1732_ NAND2
X5020 VSS VDD _1646_ _1648_ _1733_ XOR
X5021 VSS VDD _1733_ _1734_ INVERTER
X5022 VSS VDD _1247_ _1286_ _1735_ XOR
X5023 VSS VDD _1642_ _1644_ _1736_ XOR
X5024 VSS VDD _1639_ _1641_ _1737_ XOR
X5025 VSS VDD _1261_ _1279_ _1738_ XOR
X5026 VSS VDD _1737_ _1738_ _1740_ NOR2
X5027 VSS VDD _1595_ _1638_ _1741_ XOR
X5028 VSS VDD _1550_ _1633_ _1742_ NAND2
X5029 VSS VDD _1589_ _1619_ _1742_ _1743_ OAI21
X5030 VSS VDD finestra_gaussiana2_0_ sensor2_0_ _1270_ _1744_ AOI21
X5031 VSS VDD _1272_ _1589_ _1743_ _1744_ _1745_ OAI31
X5032 VSS VDD _1272_ _1589_ _1743_ _1744_ _1746_ NOR4
X5033 VSS VDD _1272_ _1274_ _1747_ XOR
X5034 VSS VDD _1745_ _1747_ _1746_ _1748_ AOI21
X5035 VSS VDD _1275_ _1278_ _1749_ XOR
X5036 VSS VDD _1741_ _1748_ _1751_ NOR2
X5037 VSS VDD _1741_ _1748_ _1749_ _1752_ AOI21
X5038 VSS VDD _1737_ _1738_ _1751_ _1752_ _1753_ AOI211
X5039 VSS VDD _1736_ _1740_ _1753_ _1754_ NOR3
X5040 VSS VDD _1740_ _1753_ _1736_ _1755_ OAI21
X5041 VSS VDD _1281_ _1282_ _1756_ XOR
X5042 VSS VDD _1755_ _1756_ _1754_ _1757_ AOI21
X5043 VSS VDD _1642_ _1643_ _1626_ _1758_ OAI21
X5044 VSS VDD _1628_ _1758_ _1759_ XOR
X5045 VSS VDD _1757_ _1759_ _1760_ NOR2
X5046 VSS VDD _1252_ _1284_ _1762_ XOR
X5047 VSS VDD _1757_ _1759_ _1762_ _1763_ AOI21
X5048 VSS VDD _1734_ _1763_ _1735_ _1760_ _1764_ OAI31
X5049 VSS VDD _1760_ _1763_ _1734_ _1765_ OAI21
X5050 VSS VDD _1764_ _1765_ _1766_ NAND2
X5051 VSS VDD _1732_ _1766_ _1731_ _1767_ AOI21
X5052 VSS VDD _1726_ _1767_ _1727_ _1768_ AOI21
X5053 VSS VDD _1723_ _1768_ _1722_ _1769_ AOI21
X5054 VSS VDD _1718_ _1769_ _1719_ _1770_ OAI21
X5055 VSS VDD _1714_ _1770_ _1771_ NOR2
X5056 VSS VDD _1713_ _1770_ _1714_ _1705_ _1773_ AOI211
X5057 VSS VDD _1704_ _1771_ _1707_ _1712_ _1774_ OAI31
X5058 VSS VDD _1698_ _1774_ _1696_ _1775_ AOI21
X5059 VSS VDD _1699_ _1704_ _1697_ _1773_ _1776_ OAI31
X5060 VSS VDD _1689_ _1776_ _1687_ _1777_ AOI21
X5061 VSS VDD _1690_ _1775_ _1688_ _1778_ OAI21
X5062 VSS VDD _1680_ _1778_ _1678_ _1779_ AOI21
X5063 VSS VDD _1681_ _1777_ _1679_ _1780_ OAI21
X5064 VSS VDD _1298_ _1305_ _1781_ XOR
X5065 VSS VDD _1298_ _1304_ _1782_ XOR
X5066 VSS VDD _1680_ _1778_ _1781_ _1678_ _1784_ AOI211
X5067 VSS VDD _1681_ _1777_ _1782_ _1679_ _1785_ OAI211
X5068 VSS VDD _1780_ _1781_ _1786_ XOR
X5069 VSS VDD _1779_ _1781_ _1787_ XOR
X5070 VSS VDD _1311_ _1787_ _1788_ NOR2
X5071 VSS VDD _1312_ _1786_ _1789_ NAND2
X5072 VSS VDD _1312_ _1785_ _1307_ _1790_ AOI21
X5073 VSS VDD _1790_ _0000__3_ INVERTER
X5074 VSS VDD _1689_ _1775_ _1791_ XOR
X5075 VSS VDD _1791_ _1792_ INVERTER
X5076 VSS VDD _1681_ _1777_ _1794_ XOR
X5077 VSS VDD _1794_ _1795_ INVERTER
X5078 VSS VDD _1780_ _1781_ _1312_ _1796_ AOI21
X5079 VSS VDD _1779_ _1782_ _1311_ _1797_ OAI21
X5080 VSS VDD _1308_ _1784_ _1798_ NOR2
X5081 VSS VDD _1307_ _1785_ _1799_ NAND2
X5082 VSS VDD _0000__3_ _1799_ _1796_ _1800_ AOI21
X5083 VSS VDD _1790_ _1798_ _1797_ _1801_ OAI21
X5084 VSS VDD _1786_ _0000__3_ _1802_ NOR2
X5085 VSS VDD _1787_ _1790_ _1803_ NAND2
X5086 VSS VDD _1788_ _1802_ _1805_ NOR2
X5087 VSS VDD _1788_ _1795_ _1802_ _1806_ NOR3
X5088 VSS VDD _1789_ _1794_ _1803_ _1807_ NAND3
X5089 VSS VDD _1789_ _1794_ _1803_ _1800_ _1808_ AOI31
X5090 VSS VDD _1808_ _0000__2_ INVERTER
X5091 VSS VDD _1795_ _1808_ _1809_ NOR2
X5092 VSS VDD _1795_ _1801_ _1810_ NAND2
X5093 VSS VDD _1795_ _1808_ _1810_ _1811_ OAI21
X5094 VSS VDD _1795_ _1808_ _1810_ _1792_ _1812_ OAI211
X5095 VSS VDD _1794_ _0000__2_ _1805_ _1813_ AOI21
X5096 VSS VDD _1805_ _1809_ _1807_ _1815_ OAI21
X5097 VSS VDD _1806_ _1813_ _1812_ _0000__1_ OAI21
X5098 VSS VDD _1812_ _1815_ _1791_ _1816_ AOI21
X5099 VSS VDD _1791_ _1806_ _1811_ _1813_ _1817_ OAI31
X5100 VSS VDD _1812_ _1817_ _1818_ NAND2
X5101 VSS VDD _1806_ _1813_ _1791_ _1819_ OAI21
X5102 VSS VDD _1698_ _1774_ _1820_ XOR
X5103 VSS VDD _1819_ _1820_ _1821_ NAND2
X5104 VSS VDD _1816_ _1821_ _1818_ _0000__0_ OAI21
X5105 VSS VDD clk _0013_ INVERTER
X5106 VSS VDD clk _0011_ INVERTER
X5107 VSS VDD clk _0009_ INVERTER
X5108 VSS VDD clk _0007_ INVERTER
X5109 VSS VDD clk _0005_ INVERTER
X5110 VSS VDD clk _0003_ INVERTER
X5111 VSS VDD clk _0001_ INVERTER
X5112 VSS VDD reset _0002_ INVERTER
X5113 VSS VDD reset _0004_ INVERTER
X5114 VSS VDD reset _0006_ INVERTER
X5115 VSS VDD reset _0008_ INVERTER
X5116 VSS VDD reset _0010_ INVERTER
X5117 VSS VDD reset _0012_ INVERTER
X5118 VSS VDD reset _0014_ INVERTER
X5119 VSS VDD _2556_ LOGIC0
X5120 VSS VDD _2557_ LOGIC0
X5121 VSS VDD _2558_ LOGIC0
X5122 VSS VDD _2559_ LOGIC0
X5123 VSS VDD _0001_ _0000__0_ central_value_0_ _0002_ DFFR
X5124 VSS VDD _0003_ _0000__1_ central_value_1_ _0004_ DFFR
X5125 VSS VDD _0005_ _0000__2_ central_value_2_ _0006_ DFFR
X5126 VSS VDD _0007_ _0000__3_ central_value_3_ _0008_ DFFR
X5127 VSS VDD _0009_ _2556_ central_value_4_ _0010_ DFFR
X5128 VSS VDD _0011_ _2557_ central_value_5_ _0012_ DFFR
X5129 VSS VDD _0013_ _2558_ central_value_6_ _0014_ DFFR
X5130 VSS VDD _0015_ _2559_ central_value_7_ _0016_ DFFR

.ENDS
